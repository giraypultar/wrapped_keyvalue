VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_keyvalue
  CLASS BLOCK ;
  FOREIGN wrapped_keyvalue ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 0.000 98.030 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 296.000 13.390 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.100 300.000 274.300 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 296.000 16.150 300.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.270 296.000 111.830 300.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 0.000 155.070 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 296.000 123.790 300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 296.000 279.270 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 0.000 91.590 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.220 4.000 127.420 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 267.660 300.000 268.860 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.340 4.000 286.540 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.190 0.000 66.750 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 296.000 158.750 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 0.000 143.110 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.030 296.000 22.590 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.740 300.000 34.940 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.900 300.000 213.100 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 0.000 285.710 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 296.000 88.830 300.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 0.000 34.550 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.500 4.000 192.700 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.900 4.000 43.100 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.510 296.000 178.070 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.060 300.000 255.260 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.980 4.000 183.180 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.910 0.000 12.470 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.780 4.000 121.980 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 75.900 300.000 77.100 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 296.000 83.310 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 296.000 29.030 300.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 0.000 114.590 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 296.000 225.910 300.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 296.000 197.390 300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 296.000 79.630 300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 290.780 300.000 291.980 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.390 296.000 259.950 300.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.860 4.000 160.060 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 296.000 237.870 300.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.420 300.000 222.620 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.660 4.000 234.860 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.660 300.000 132.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.230 0.000 31.790 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 0.000 266.390 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.190 296.000 66.750 300.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.940 4.000 164.140 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 66.380 300.000 67.580 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.580 4.000 60.780 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 296.000 145.870 300.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 296.000 114.590 300.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.790 0.000 117.350 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.820 4.000 5.020 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 0.000 86.070 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.950 0.000 253.510 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.060 4.000 187.260 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.220 300.000 161.420 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 0.000 291.230 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 0.000 224.990 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.140 4.000 89.340 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.260 300.000 180.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 0.000 69.510 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.790 296.000 117.350 300.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 296.000 257.190 300.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 183.340 300.000 184.540 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 0.000 139.430 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 0.000 294.910 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 0.000 60.310 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.300 300.000 63.500 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 296.000 143.110 300.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.700 4.000 253.900 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.860 4.000 24.060 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 296.000 152.310 300.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.030 0.000 275.590 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.620 300.000 147.820 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 0.000 79.630 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.950 296.000 92.510 300.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 0.000 228.670 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.420 4.000 290.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.780 300.000 155.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 296.220 300.000 297.420 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.990 296.000 149.550 300.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.980 300.000 217.180 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.990 296.000 241.550 300.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.590 296.000 292.150 300.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 296.000 98.950 300.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.780 300.000 53.980 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 296.000 209.350 300.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 296.000 294.910 300.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.390 0.000 259.950 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 56.860 300.000 58.060 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 0.000 209.350 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.230 296.000 54.790 300.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 0.000 183.590 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.030 0.000 22.590 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 296.000 26.270 300.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.460 300.000 105.660 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 0.000 63.070 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 0.000 244.310 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.580 4.000 196.780 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.860 4.000 296.060 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 296.000 174.390 300.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 296.000 219.470 300.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 0.000 47.430 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.540 300.000 245.740 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 296.000 180.830 300.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 0.000 177.150 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 0.000 200.150 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.350 0.000 110.910 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 296.000 202.910 300.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.300 300.000 165.500 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.820 300.000 39.020 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.830 296.000 105.390 300.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 296.000 35.470 300.000 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 296.000 51.110 300.000 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.220 4.000 229.420 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.620 4.000 79.820 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.980 4.000 47.180 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 202.380 300.000 203.580 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 0.000 16.150 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.150 0.000 101.710 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 296.000 285.710 300.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 296.000 121.030 300.000 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 0.000 231.430 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 296.000 95.270 300.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.380 4.000 33.580 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.420 300.000 86.620 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.300 4.000 267.500 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.260 300.000 282.460 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 296.000 3.270 300.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 0.000 205.670 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 0.000 247.070 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.180 300.000 142.380 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 296.000 162.430 300.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 0.000 288.470 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 0.000 269.150 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 296.000 165.190 300.000 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.620 300.000 11.820 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.060 4.000 51.260 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 14.700 300.000 15.900 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 296.000 38.230 300.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.260 4.000 112.460 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 0.000 44.670 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 0.000 158.750 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 296.000 247.990 300.000 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.910 296.000 127.470 300.000 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.820 300.000 175.020 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.100 4.000 70.300 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 230.940 300.000 232.140 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.430 296.000 155.990 300.000 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.220 4.000 93.420 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 296.000 44.670 300.000 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 296.000 86.070 300.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.820 4.000 277.020 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.700 300.000 151.900 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.740 300.000 170.940 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.380 4.000 271.580 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.510 296.000 270.070 300.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.620 300.000 113.820 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 0.000 104.470 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 296.000 19.830 300.000 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 296.000 235.110 300.000 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.300 4.000 131.500 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.460 4.000 37.660 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.590 0.000 108.150 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 0.000 218.550 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.860 300.000 194.060 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 0.000 237.870 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.820 4.000 141.020 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 0.000 6.030 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 0.000 40.990 4.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.500 4.000 56.700 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.950 296.000 184.510 300.000 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 0.000 171.630 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 0.000 82.390 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 0.000 161.510 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.300 300.000 29.500 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 296.000 0.510 300.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 0.000 167.950 4.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.670 296.000 222.230 300.000 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 0.000 215.790 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.980 300.000 81.180 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 296.000 298.590 300.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 43.260 300.000 44.460 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.620 4.000 215.820 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.100 300.000 240.300 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.070 0.000 240.630 4.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.270 296.000 272.830 300.000 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 0.000 202.910 4.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 296.000 193.710 300.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 0.000 29.030 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 296.000 9.710 300.000 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 0.000 123.790 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 296.000 60.310 300.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.990 0.000 57.550 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 0.000 212.110 4.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 296.000 200.150 300.000 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.580 300.000 264.780 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.590 296.000 108.150 300.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.430 296.000 63.990 300.000 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 296.000 206.590 300.000 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.150 0.000 262.710 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 296.000 168.870 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.180 300.000 6.380 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 296.000 276.510 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 296.000 228.670 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 296.000 73.190 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.870 296.000 70.430 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.100 300.000 138.300 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.060 300.000 119.260 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 0.000 145.870 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.940 300.000 96.140 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.670 0.000 222.230 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.070 296.000 263.630 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.140 300.000 259.340 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.670 0.000 130.230 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 0.000 187.270 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.470 0.000 282.030 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 296.000 136.670 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 0.000 126.550 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 0.000 25.350 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 296.000 187.270 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.020 300.000 100.220 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.500 300.000 226.700 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 0.000 88.830 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 296.000 288.470 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.340 300.000 48.540 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.420 4.000 18.620 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.180 4.000 244.380 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 0.000 174.390 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 0.000 73.190 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.630 0.000 234.190 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 0.000 297.670 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 296.000 171.630 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.020 4.000 66.220 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 296.000 41.910 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.990 296.000 57.550 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 296.000 48.350 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.740 4.000 102.940 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.500 300.000 90.700 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 0.000 136.670 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 296.000 250.750 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 286.700 300.000 287.900 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.150 296.000 101.710 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.100 4.000 206.300 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.460 4.000 173.660 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.180 300.000 278.380 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.900 4.000 281.100 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.780 300.000 189.980 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.180 4.000 108.380 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.390 296.000 282.950 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 296.000 140.350 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.390 0.000 75.950 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.580 300.000 128.780 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.910 0.000 196.470 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.140 300.000 21.340 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.260 4.000 248.460 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 0.000 250.750 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 0.000 38.230 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 0.000 120.110 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.460 300.000 71.660 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 296.000 266.390 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.020 300.000 236.220 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 0.000 257.190 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.660 4.000 98.860 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.140 300.000 123.340 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 0.000 3.270 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.620 300.000 249.820 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.870 296.000 254.430 300.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.270 0.000 272.830 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 296.000 244.310 300.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.380 4.000 135.580 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 0.000 165.190 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 0.000 193.710 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.670 296.000 130.230 300.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.900 4.000 145.100 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 0.000 51.110 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 296.000 190.950 300.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 296.000 133.910 300.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 0.000 132.990 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 296.000 231.430 300.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 24.220 300.000 25.420 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.780 4.000 257.980 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 206.460 300.000 207.660 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 0.000 53.870 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 0.000 95.270 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 0.000 148.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 196.940 300.000 198.140 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 0.000 152.310 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 296.000 215.790 300.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 296.000 213.030 300.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.230 296.000 31.790 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 296.000 76.870 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 0.000 180.830 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.060 4.000 85.260 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 296.000 6.950 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.540 300.000 109.740 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 4.285 4.845 299.775 290.615 ;
      LAYER met1 ;
        RECT 0.070 0.380 299.850 298.480 ;
      LAYER met2 ;
        RECT 0.790 295.720 2.430 298.510 ;
        RECT 3.550 295.720 6.110 298.510 ;
        RECT 7.230 295.720 8.870 298.510 ;
        RECT 9.990 295.720 12.550 298.510 ;
        RECT 13.670 295.720 15.310 298.510 ;
        RECT 16.430 295.720 18.990 298.510 ;
        RECT 20.110 295.720 21.750 298.510 ;
        RECT 22.870 295.720 25.430 298.510 ;
        RECT 26.550 295.720 28.190 298.510 ;
        RECT 29.310 295.720 30.950 298.510 ;
        RECT 32.070 295.720 34.630 298.510 ;
        RECT 35.750 295.720 37.390 298.510 ;
        RECT 38.510 295.720 41.070 298.510 ;
        RECT 42.190 295.720 43.830 298.510 ;
        RECT 44.950 295.720 47.510 298.510 ;
        RECT 48.630 295.720 50.270 298.510 ;
        RECT 51.390 295.720 53.950 298.510 ;
        RECT 55.070 295.720 56.710 298.510 ;
        RECT 57.830 295.720 59.470 298.510 ;
        RECT 60.590 295.720 63.150 298.510 ;
        RECT 64.270 295.720 65.910 298.510 ;
        RECT 67.030 295.720 69.590 298.510 ;
        RECT 70.710 295.720 72.350 298.510 ;
        RECT 73.470 295.720 76.030 298.510 ;
        RECT 77.150 295.720 78.790 298.510 ;
        RECT 79.910 295.720 82.470 298.510 ;
        RECT 83.590 295.720 85.230 298.510 ;
        RECT 86.350 295.720 87.990 298.510 ;
        RECT 89.110 295.720 91.670 298.510 ;
        RECT 92.790 295.720 94.430 298.510 ;
        RECT 95.550 295.720 98.110 298.510 ;
        RECT 99.230 295.720 100.870 298.510 ;
        RECT 101.990 295.720 104.550 298.510 ;
        RECT 105.670 295.720 107.310 298.510 ;
        RECT 108.430 295.720 110.990 298.510 ;
        RECT 112.110 295.720 113.750 298.510 ;
        RECT 114.870 295.720 116.510 298.510 ;
        RECT 117.630 295.720 120.190 298.510 ;
        RECT 121.310 295.720 122.950 298.510 ;
        RECT 124.070 295.720 126.630 298.510 ;
        RECT 127.750 295.720 129.390 298.510 ;
        RECT 130.510 295.720 133.070 298.510 ;
        RECT 134.190 295.720 135.830 298.510 ;
        RECT 136.950 295.720 139.510 298.510 ;
        RECT 140.630 295.720 142.270 298.510 ;
        RECT 143.390 295.720 145.030 298.510 ;
        RECT 146.150 295.720 148.710 298.510 ;
        RECT 149.830 295.720 151.470 298.510 ;
        RECT 152.590 295.720 155.150 298.510 ;
        RECT 156.270 295.720 157.910 298.510 ;
        RECT 159.030 295.720 161.590 298.510 ;
        RECT 162.710 295.720 164.350 298.510 ;
        RECT 165.470 295.720 168.030 298.510 ;
        RECT 169.150 295.720 170.790 298.510 ;
        RECT 171.910 295.720 173.550 298.510 ;
        RECT 174.670 295.720 177.230 298.510 ;
        RECT 178.350 295.720 179.990 298.510 ;
        RECT 181.110 295.720 183.670 298.510 ;
        RECT 184.790 295.720 186.430 298.510 ;
        RECT 187.550 295.720 190.110 298.510 ;
        RECT 191.230 295.720 192.870 298.510 ;
        RECT 193.990 295.720 196.550 298.510 ;
        RECT 197.670 295.720 199.310 298.510 ;
        RECT 200.430 295.720 202.070 298.510 ;
        RECT 203.190 295.720 205.750 298.510 ;
        RECT 206.870 295.720 208.510 298.510 ;
        RECT 209.630 295.720 212.190 298.510 ;
        RECT 213.310 295.720 214.950 298.510 ;
        RECT 216.070 295.720 218.630 298.510 ;
        RECT 219.750 295.720 221.390 298.510 ;
        RECT 222.510 295.720 225.070 298.510 ;
        RECT 226.190 295.720 227.830 298.510 ;
        RECT 228.950 295.720 230.590 298.510 ;
        RECT 231.710 295.720 234.270 298.510 ;
        RECT 235.390 295.720 237.030 298.510 ;
        RECT 238.150 295.720 240.710 298.510 ;
        RECT 241.830 295.720 243.470 298.510 ;
        RECT 244.590 295.720 247.150 298.510 ;
        RECT 248.270 295.720 249.910 298.510 ;
        RECT 251.030 295.720 253.590 298.510 ;
        RECT 254.710 295.720 256.350 298.510 ;
        RECT 257.470 295.720 259.110 298.510 ;
        RECT 260.230 295.720 262.790 298.510 ;
        RECT 263.910 295.720 265.550 298.510 ;
        RECT 266.670 295.720 269.230 298.510 ;
        RECT 270.350 295.720 271.990 298.510 ;
        RECT 273.110 295.720 275.670 298.510 ;
        RECT 276.790 295.720 278.430 298.510 ;
        RECT 279.550 295.720 282.110 298.510 ;
        RECT 283.230 295.720 284.870 298.510 ;
        RECT 285.990 295.720 287.630 298.510 ;
        RECT 288.750 295.720 291.310 298.510 ;
        RECT 292.430 295.720 294.070 298.510 ;
        RECT 295.190 295.720 297.750 298.510 ;
        RECT 298.870 295.720 299.820 298.510 ;
        RECT 0.090 4.280 299.820 295.720 ;
        RECT 0.790 0.155 2.430 4.280 ;
        RECT 3.550 0.155 5.190 4.280 ;
        RECT 6.310 0.155 8.870 4.280 ;
        RECT 9.990 0.155 11.630 4.280 ;
        RECT 12.750 0.155 15.310 4.280 ;
        RECT 16.430 0.155 18.070 4.280 ;
        RECT 19.190 0.155 21.750 4.280 ;
        RECT 22.870 0.155 24.510 4.280 ;
        RECT 25.630 0.155 28.190 4.280 ;
        RECT 29.310 0.155 30.950 4.280 ;
        RECT 32.070 0.155 33.710 4.280 ;
        RECT 34.830 0.155 37.390 4.280 ;
        RECT 38.510 0.155 40.150 4.280 ;
        RECT 41.270 0.155 43.830 4.280 ;
        RECT 44.950 0.155 46.590 4.280 ;
        RECT 47.710 0.155 50.270 4.280 ;
        RECT 51.390 0.155 53.030 4.280 ;
        RECT 54.150 0.155 56.710 4.280 ;
        RECT 57.830 0.155 59.470 4.280 ;
        RECT 60.590 0.155 62.230 4.280 ;
        RECT 63.350 0.155 65.910 4.280 ;
        RECT 67.030 0.155 68.670 4.280 ;
        RECT 69.790 0.155 72.350 4.280 ;
        RECT 73.470 0.155 75.110 4.280 ;
        RECT 76.230 0.155 78.790 4.280 ;
        RECT 79.910 0.155 81.550 4.280 ;
        RECT 82.670 0.155 85.230 4.280 ;
        RECT 86.350 0.155 87.990 4.280 ;
        RECT 89.110 0.155 90.750 4.280 ;
        RECT 91.870 0.155 94.430 4.280 ;
        RECT 95.550 0.155 97.190 4.280 ;
        RECT 98.310 0.155 100.870 4.280 ;
        RECT 101.990 0.155 103.630 4.280 ;
        RECT 104.750 0.155 107.310 4.280 ;
        RECT 108.430 0.155 110.070 4.280 ;
        RECT 111.190 0.155 113.750 4.280 ;
        RECT 114.870 0.155 116.510 4.280 ;
        RECT 117.630 0.155 119.270 4.280 ;
        RECT 120.390 0.155 122.950 4.280 ;
        RECT 124.070 0.155 125.710 4.280 ;
        RECT 126.830 0.155 129.390 4.280 ;
        RECT 130.510 0.155 132.150 4.280 ;
        RECT 133.270 0.155 135.830 4.280 ;
        RECT 136.950 0.155 138.590 4.280 ;
        RECT 139.710 0.155 142.270 4.280 ;
        RECT 143.390 0.155 145.030 4.280 ;
        RECT 146.150 0.155 147.790 4.280 ;
        RECT 148.910 0.155 151.470 4.280 ;
        RECT 152.590 0.155 154.230 4.280 ;
        RECT 155.350 0.155 157.910 4.280 ;
        RECT 159.030 0.155 160.670 4.280 ;
        RECT 161.790 0.155 164.350 4.280 ;
        RECT 165.470 0.155 167.110 4.280 ;
        RECT 168.230 0.155 170.790 4.280 ;
        RECT 171.910 0.155 173.550 4.280 ;
        RECT 174.670 0.155 176.310 4.280 ;
        RECT 177.430 0.155 179.990 4.280 ;
        RECT 181.110 0.155 182.750 4.280 ;
        RECT 183.870 0.155 186.430 4.280 ;
        RECT 187.550 0.155 189.190 4.280 ;
        RECT 190.310 0.155 192.870 4.280 ;
        RECT 193.990 0.155 195.630 4.280 ;
        RECT 196.750 0.155 199.310 4.280 ;
        RECT 200.430 0.155 202.070 4.280 ;
        RECT 203.190 0.155 204.830 4.280 ;
        RECT 205.950 0.155 208.510 4.280 ;
        RECT 209.630 0.155 211.270 4.280 ;
        RECT 212.390 0.155 214.950 4.280 ;
        RECT 216.070 0.155 217.710 4.280 ;
        RECT 218.830 0.155 221.390 4.280 ;
        RECT 222.510 0.155 224.150 4.280 ;
        RECT 225.270 0.155 227.830 4.280 ;
        RECT 228.950 0.155 230.590 4.280 ;
        RECT 231.710 0.155 233.350 4.280 ;
        RECT 234.470 0.155 237.030 4.280 ;
        RECT 238.150 0.155 239.790 4.280 ;
        RECT 240.910 0.155 243.470 4.280 ;
        RECT 244.590 0.155 246.230 4.280 ;
        RECT 247.350 0.155 249.910 4.280 ;
        RECT 251.030 0.155 252.670 4.280 ;
        RECT 253.790 0.155 256.350 4.280 ;
        RECT 257.470 0.155 259.110 4.280 ;
        RECT 260.230 0.155 261.870 4.280 ;
        RECT 262.990 0.155 265.550 4.280 ;
        RECT 266.670 0.155 268.310 4.280 ;
        RECT 269.430 0.155 271.990 4.280 ;
        RECT 273.110 0.155 274.750 4.280 ;
        RECT 275.870 0.155 278.430 4.280 ;
        RECT 279.550 0.155 281.190 4.280 ;
        RECT 282.310 0.155 284.870 4.280 ;
        RECT 285.990 0.155 287.630 4.280 ;
        RECT 288.750 0.155 290.390 4.280 ;
        RECT 291.510 0.155 294.070 4.280 ;
        RECT 295.190 0.155 296.830 4.280 ;
        RECT 297.950 0.155 299.820 4.280 ;
      LAYER met3 ;
        RECT 0.065 296.460 295.600 296.985 ;
        RECT 4.400 295.820 295.600 296.460 ;
        RECT 4.400 294.460 296.635 295.820 ;
        RECT 0.065 292.380 296.635 294.460 ;
        RECT 0.065 291.020 295.600 292.380 ;
        RECT 4.400 290.380 295.600 291.020 ;
        RECT 4.400 289.020 296.635 290.380 ;
        RECT 0.065 288.300 296.635 289.020 ;
        RECT 0.065 286.940 295.600 288.300 ;
        RECT 4.400 286.300 295.600 286.940 ;
        RECT 4.400 284.940 296.635 286.300 ;
        RECT 0.065 282.860 296.635 284.940 ;
        RECT 0.065 281.500 295.600 282.860 ;
        RECT 4.400 280.860 295.600 281.500 ;
        RECT 4.400 279.500 296.635 280.860 ;
        RECT 0.065 278.780 296.635 279.500 ;
        RECT 0.065 277.420 295.600 278.780 ;
        RECT 4.400 276.780 295.600 277.420 ;
        RECT 4.400 275.420 296.635 276.780 ;
        RECT 0.065 274.700 296.635 275.420 ;
        RECT 0.065 272.700 295.600 274.700 ;
        RECT 0.065 271.980 296.635 272.700 ;
        RECT 4.400 269.980 296.635 271.980 ;
        RECT 0.065 269.260 296.635 269.980 ;
        RECT 0.065 267.900 295.600 269.260 ;
        RECT 4.400 267.260 295.600 267.900 ;
        RECT 4.400 265.900 296.635 267.260 ;
        RECT 0.065 265.180 296.635 265.900 ;
        RECT 0.065 263.180 295.600 265.180 ;
        RECT 0.065 262.460 296.635 263.180 ;
        RECT 4.400 260.460 296.635 262.460 ;
        RECT 0.065 259.740 296.635 260.460 ;
        RECT 0.065 258.380 295.600 259.740 ;
        RECT 4.400 257.740 295.600 258.380 ;
        RECT 4.400 256.380 296.635 257.740 ;
        RECT 0.065 255.660 296.635 256.380 ;
        RECT 0.065 254.300 295.600 255.660 ;
        RECT 4.400 253.660 295.600 254.300 ;
        RECT 4.400 252.300 296.635 253.660 ;
        RECT 0.065 250.220 296.635 252.300 ;
        RECT 0.065 248.860 295.600 250.220 ;
        RECT 4.400 248.220 295.600 248.860 ;
        RECT 4.400 246.860 296.635 248.220 ;
        RECT 0.065 246.140 296.635 246.860 ;
        RECT 0.065 244.780 295.600 246.140 ;
        RECT 4.400 244.140 295.600 244.780 ;
        RECT 4.400 242.780 296.635 244.140 ;
        RECT 0.065 240.700 296.635 242.780 ;
        RECT 0.065 239.340 295.600 240.700 ;
        RECT 4.400 238.700 295.600 239.340 ;
        RECT 4.400 237.340 296.635 238.700 ;
        RECT 0.065 236.620 296.635 237.340 ;
        RECT 0.065 235.260 295.600 236.620 ;
        RECT 4.400 234.620 295.600 235.260 ;
        RECT 4.400 233.260 296.635 234.620 ;
        RECT 0.065 232.540 296.635 233.260 ;
        RECT 0.065 230.540 295.600 232.540 ;
        RECT 0.065 229.820 296.635 230.540 ;
        RECT 4.400 227.820 296.635 229.820 ;
        RECT 0.065 227.100 296.635 227.820 ;
        RECT 0.065 225.740 295.600 227.100 ;
        RECT 4.400 225.100 295.600 225.740 ;
        RECT 4.400 223.740 296.635 225.100 ;
        RECT 0.065 223.020 296.635 223.740 ;
        RECT 0.065 221.020 295.600 223.020 ;
        RECT 0.065 220.300 296.635 221.020 ;
        RECT 4.400 218.300 296.635 220.300 ;
        RECT 0.065 217.580 296.635 218.300 ;
        RECT 0.065 216.220 295.600 217.580 ;
        RECT 4.400 215.580 295.600 216.220 ;
        RECT 4.400 214.220 296.635 215.580 ;
        RECT 0.065 213.500 296.635 214.220 ;
        RECT 0.065 212.140 295.600 213.500 ;
        RECT 4.400 211.500 295.600 212.140 ;
        RECT 4.400 210.140 296.635 211.500 ;
        RECT 0.065 208.060 296.635 210.140 ;
        RECT 0.065 206.700 295.600 208.060 ;
        RECT 4.400 206.060 295.600 206.700 ;
        RECT 4.400 204.700 296.635 206.060 ;
        RECT 0.065 203.980 296.635 204.700 ;
        RECT 0.065 202.620 295.600 203.980 ;
        RECT 4.400 201.980 295.600 202.620 ;
        RECT 4.400 200.620 296.635 201.980 ;
        RECT 0.065 198.540 296.635 200.620 ;
        RECT 0.065 197.180 295.600 198.540 ;
        RECT 4.400 196.540 295.600 197.180 ;
        RECT 4.400 195.180 296.635 196.540 ;
        RECT 0.065 194.460 296.635 195.180 ;
        RECT 0.065 193.100 295.600 194.460 ;
        RECT 4.400 192.460 295.600 193.100 ;
        RECT 4.400 191.100 296.635 192.460 ;
        RECT 0.065 190.380 296.635 191.100 ;
        RECT 0.065 188.380 295.600 190.380 ;
        RECT 0.065 187.660 296.635 188.380 ;
        RECT 4.400 185.660 296.635 187.660 ;
        RECT 0.065 184.940 296.635 185.660 ;
        RECT 0.065 183.580 295.600 184.940 ;
        RECT 4.400 182.940 295.600 183.580 ;
        RECT 4.400 181.580 296.635 182.940 ;
        RECT 0.065 180.860 296.635 181.580 ;
        RECT 0.065 178.860 295.600 180.860 ;
        RECT 0.065 178.140 296.635 178.860 ;
        RECT 4.400 176.140 296.635 178.140 ;
        RECT 0.065 175.420 296.635 176.140 ;
        RECT 0.065 174.060 295.600 175.420 ;
        RECT 4.400 173.420 295.600 174.060 ;
        RECT 4.400 172.060 296.635 173.420 ;
        RECT 0.065 171.340 296.635 172.060 ;
        RECT 0.065 169.980 295.600 171.340 ;
        RECT 4.400 169.340 295.600 169.980 ;
        RECT 4.400 167.980 296.635 169.340 ;
        RECT 0.065 165.900 296.635 167.980 ;
        RECT 0.065 164.540 295.600 165.900 ;
        RECT 4.400 163.900 295.600 164.540 ;
        RECT 4.400 162.540 296.635 163.900 ;
        RECT 0.065 161.820 296.635 162.540 ;
        RECT 0.065 160.460 295.600 161.820 ;
        RECT 4.400 159.820 295.600 160.460 ;
        RECT 4.400 158.460 296.635 159.820 ;
        RECT 0.065 156.380 296.635 158.460 ;
        RECT 0.065 155.020 295.600 156.380 ;
        RECT 4.400 154.380 295.600 155.020 ;
        RECT 4.400 153.020 296.635 154.380 ;
        RECT 0.065 152.300 296.635 153.020 ;
        RECT 0.065 150.940 295.600 152.300 ;
        RECT 4.400 150.300 295.600 150.940 ;
        RECT 4.400 148.940 296.635 150.300 ;
        RECT 0.065 148.220 296.635 148.940 ;
        RECT 0.065 146.220 295.600 148.220 ;
        RECT 0.065 145.500 296.635 146.220 ;
        RECT 4.400 143.500 296.635 145.500 ;
        RECT 0.065 142.780 296.635 143.500 ;
        RECT 0.065 141.420 295.600 142.780 ;
        RECT 4.400 140.780 295.600 141.420 ;
        RECT 4.400 139.420 296.635 140.780 ;
        RECT 0.065 138.700 296.635 139.420 ;
        RECT 0.065 136.700 295.600 138.700 ;
        RECT 0.065 135.980 296.635 136.700 ;
        RECT 4.400 133.980 296.635 135.980 ;
        RECT 0.065 133.260 296.635 133.980 ;
        RECT 0.065 131.900 295.600 133.260 ;
        RECT 4.400 131.260 295.600 131.900 ;
        RECT 4.400 129.900 296.635 131.260 ;
        RECT 0.065 129.180 296.635 129.900 ;
        RECT 0.065 127.820 295.600 129.180 ;
        RECT 4.400 127.180 295.600 127.820 ;
        RECT 4.400 125.820 296.635 127.180 ;
        RECT 0.065 123.740 296.635 125.820 ;
        RECT 0.065 122.380 295.600 123.740 ;
        RECT 4.400 121.740 295.600 122.380 ;
        RECT 4.400 120.380 296.635 121.740 ;
        RECT 0.065 119.660 296.635 120.380 ;
        RECT 0.065 118.300 295.600 119.660 ;
        RECT 4.400 117.660 295.600 118.300 ;
        RECT 4.400 116.300 296.635 117.660 ;
        RECT 0.065 114.220 296.635 116.300 ;
        RECT 0.065 112.860 295.600 114.220 ;
        RECT 4.400 112.220 295.600 112.860 ;
        RECT 4.400 110.860 296.635 112.220 ;
        RECT 0.065 110.140 296.635 110.860 ;
        RECT 0.065 108.780 295.600 110.140 ;
        RECT 4.400 108.140 295.600 108.780 ;
        RECT 4.400 106.780 296.635 108.140 ;
        RECT 0.065 106.060 296.635 106.780 ;
        RECT 0.065 104.060 295.600 106.060 ;
        RECT 0.065 103.340 296.635 104.060 ;
        RECT 4.400 101.340 296.635 103.340 ;
        RECT 0.065 100.620 296.635 101.340 ;
        RECT 0.065 99.260 295.600 100.620 ;
        RECT 4.400 98.620 295.600 99.260 ;
        RECT 4.400 97.260 296.635 98.620 ;
        RECT 0.065 96.540 296.635 97.260 ;
        RECT 0.065 94.540 295.600 96.540 ;
        RECT 0.065 93.820 296.635 94.540 ;
        RECT 4.400 91.820 296.635 93.820 ;
        RECT 0.065 91.100 296.635 91.820 ;
        RECT 0.065 89.740 295.600 91.100 ;
        RECT 4.400 89.100 295.600 89.740 ;
        RECT 4.400 87.740 296.635 89.100 ;
        RECT 0.065 87.020 296.635 87.740 ;
        RECT 0.065 85.660 295.600 87.020 ;
        RECT 4.400 85.020 295.600 85.660 ;
        RECT 4.400 83.660 296.635 85.020 ;
        RECT 0.065 81.580 296.635 83.660 ;
        RECT 0.065 80.220 295.600 81.580 ;
        RECT 4.400 79.580 295.600 80.220 ;
        RECT 4.400 78.220 296.635 79.580 ;
        RECT 0.065 77.500 296.635 78.220 ;
        RECT 0.065 76.140 295.600 77.500 ;
        RECT 4.400 75.500 295.600 76.140 ;
        RECT 4.400 74.140 296.635 75.500 ;
        RECT 0.065 72.060 296.635 74.140 ;
        RECT 0.065 70.700 295.600 72.060 ;
        RECT 4.400 70.060 295.600 70.700 ;
        RECT 4.400 68.700 296.635 70.060 ;
        RECT 0.065 67.980 296.635 68.700 ;
        RECT 0.065 66.620 295.600 67.980 ;
        RECT 4.400 65.980 295.600 66.620 ;
        RECT 4.400 64.620 296.635 65.980 ;
        RECT 0.065 63.900 296.635 64.620 ;
        RECT 0.065 61.900 295.600 63.900 ;
        RECT 0.065 61.180 296.635 61.900 ;
        RECT 4.400 59.180 296.635 61.180 ;
        RECT 0.065 58.460 296.635 59.180 ;
        RECT 0.065 57.100 295.600 58.460 ;
        RECT 4.400 56.460 295.600 57.100 ;
        RECT 4.400 55.100 296.635 56.460 ;
        RECT 0.065 54.380 296.635 55.100 ;
        RECT 0.065 52.380 295.600 54.380 ;
        RECT 0.065 51.660 296.635 52.380 ;
        RECT 4.400 49.660 296.635 51.660 ;
        RECT 0.065 48.940 296.635 49.660 ;
        RECT 0.065 47.580 295.600 48.940 ;
        RECT 4.400 46.940 295.600 47.580 ;
        RECT 4.400 45.580 296.635 46.940 ;
        RECT 0.065 44.860 296.635 45.580 ;
        RECT 0.065 43.500 295.600 44.860 ;
        RECT 4.400 42.860 295.600 43.500 ;
        RECT 4.400 41.500 296.635 42.860 ;
        RECT 0.065 39.420 296.635 41.500 ;
        RECT 0.065 38.060 295.600 39.420 ;
        RECT 4.400 37.420 295.600 38.060 ;
        RECT 4.400 36.060 296.635 37.420 ;
        RECT 0.065 35.340 296.635 36.060 ;
        RECT 0.065 33.980 295.600 35.340 ;
        RECT 4.400 33.340 295.600 33.980 ;
        RECT 4.400 31.980 296.635 33.340 ;
        RECT 0.065 29.900 296.635 31.980 ;
        RECT 0.065 28.540 295.600 29.900 ;
        RECT 4.400 27.900 295.600 28.540 ;
        RECT 4.400 26.540 296.635 27.900 ;
        RECT 0.065 25.820 296.635 26.540 ;
        RECT 0.065 24.460 295.600 25.820 ;
        RECT 4.400 23.820 295.600 24.460 ;
        RECT 4.400 22.460 296.635 23.820 ;
        RECT 0.065 21.740 296.635 22.460 ;
        RECT 0.065 19.740 295.600 21.740 ;
        RECT 0.065 19.020 296.635 19.740 ;
        RECT 4.400 17.020 296.635 19.020 ;
        RECT 0.065 16.300 296.635 17.020 ;
        RECT 0.065 14.940 295.600 16.300 ;
        RECT 4.400 14.300 295.600 14.940 ;
        RECT 4.400 12.940 296.635 14.300 ;
        RECT 0.065 12.220 296.635 12.940 ;
        RECT 0.065 10.220 295.600 12.220 ;
        RECT 0.065 9.500 296.635 10.220 ;
        RECT 4.400 7.500 296.635 9.500 ;
        RECT 0.065 6.780 296.635 7.500 ;
        RECT 0.065 5.420 295.600 6.780 ;
        RECT 4.400 4.780 295.600 5.420 ;
        RECT 4.400 3.420 296.635 4.780 ;
        RECT 0.065 2.700 296.635 3.420 ;
        RECT 0.065 0.700 295.600 2.700 ;
        RECT 0.065 0.175 296.635 0.700 ;
      LAYER met4 ;
        RECT 0.295 288.960 295.025 294.265 ;
        RECT 0.295 10.240 20.640 288.960 ;
        RECT 23.040 10.240 97.440 288.960 ;
        RECT 99.840 10.240 174.240 288.960 ;
        RECT 176.640 10.240 251.040 288.960 ;
        RECT 253.440 10.240 295.025 288.960 ;
        RECT 0.295 0.855 295.025 10.240 ;
  END
END wrapped_keyvalue
END LIBRARY

