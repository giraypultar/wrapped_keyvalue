/* Machine-generated using Migen */
module keyvalue_3(
	input [63:0] KEY_i,
	input [63:0] VALUE_i_o,
	input [3:0] SEL_i,
	input [63:0] ADR_i,
	input [63:0] DAT_i,
	input WE_i,
	input STB_i,
	input CYC_i,
	output reg STALL_o,
	output reg ACK_o,
	output reg [63:0] DAT_o,
	output [63:0] LA_o,
	input sys_clk,
	input sys_rst
);

reg [63:0] storak0 = 64'd0;
reg [63:0] storak1 = 64'd0;
reg [63:0] storak2 = 64'd0;
reg [63:0] storak3 = 64'd0;
reg [63:0] storak4 = 64'd0;
reg [63:0] storak5 = 64'd0;
reg [63:0] storak6 = 64'd0;
reg [63:0] storak7 = 64'd0;
reg [63:0] storak8 = 64'd0;
reg [63:0] storak9 = 64'd0;
reg [63:0] storak10 = 64'd0;
reg [63:0] storak11 = 64'd0;
reg [63:0] storak12 = 64'd0;
reg [63:0] storak13 = 64'd0;
reg [63:0] storak14 = 64'd0;
reg [63:0] storak15 = 64'd0;
reg [63:0] storak16 = 64'd0;
reg [63:0] storak17 = 64'd0;
reg [63:0] storak18 = 64'd0;
reg [63:0] storak19 = 64'd0;
reg [63:0] storak20 = 64'd0;
reg [63:0] storak21 = 64'd0;
reg [63:0] storak22 = 64'd0;
reg [63:0] storak23 = 64'd0;
reg [63:0] storak24 = 64'd0;
reg [63:0] storak25 = 64'd0;
reg [63:0] storak26 = 64'd0;
reg [63:0] storak27 = 64'd0;
reg [63:0] storak28 = 64'd0;
reg [63:0] storak29 = 64'd0;
reg [63:0] storak30 = 64'd0;
reg [63:0] storak31 = 64'd0;
reg [63:0] storak32 = 64'd0;
reg [63:0] storak33 = 64'd0;
reg [63:0] storak34 = 64'd0;
reg [63:0] storak35 = 64'd0;
reg [63:0] storak36 = 64'd0;
reg [63:0] storak37 = 64'd0;
reg [63:0] storak38 = 64'd0;
reg [63:0] storak39 = 64'd0;
reg [63:0] storak40 = 64'd0;
reg [63:0] storak41 = 64'd0;
reg [63:0] storak42 = 64'd0;
reg [63:0] storak43 = 64'd0;
reg [63:0] storak44 = 64'd0;
reg [63:0] storak45 = 64'd0;
reg [63:0] storak46 = 64'd0;
reg [63:0] storak47 = 64'd0;
reg [63:0] storak48 = 64'd0;
reg [63:0] storak49 = 64'd0;
reg [63:0] storak50 = 64'd0;
reg [63:0] storak51 = 64'd0;
reg [63:0] storak52 = 64'd0;
reg [63:0] storak53 = 64'd0;
reg [63:0] storak54 = 64'd0;
reg [63:0] storak55 = 64'd0;
reg [63:0] storak56 = 64'd0;
reg [63:0] storak57 = 64'd0;
reg [63:0] storak58 = 64'd0;
reg [63:0] storak59 = 64'd0;
reg [63:0] storak60 = 64'd0;
reg [63:0] storak61 = 64'd0;
reg [63:0] storak62 = 64'd0;
reg [63:0] storak63 = 64'd0;
reg [63:0] storak64 = 64'd0;
reg [63:0] storak65 = 64'd0;
reg [63:0] storak66 = 64'd0;
reg [63:0] storak67 = 64'd0;
reg [63:0] storak68 = 64'd0;
reg [63:0] storak69 = 64'd0;
reg [63:0] storak70 = 64'd0;
reg [63:0] storak71 = 64'd0;
reg [63:0] storak72 = 64'd0;
reg [63:0] storak73 = 64'd0;
reg [63:0] storak74 = 64'd0;
reg [63:0] storak75 = 64'd0;
reg [63:0] storak76 = 64'd0;
reg [63:0] storak77 = 64'd0;
reg [63:0] storak78 = 64'd0;
reg [63:0] storak79 = 64'd0;
reg [63:0] storak80 = 64'd0;
reg [63:0] storak81 = 64'd0;
reg [63:0] storak82 = 64'd0;
reg [63:0] storak83 = 64'd0;
reg [63:0] storak84 = 64'd0;
reg [63:0] storak85 = 64'd0;
reg [63:0] storak86 = 64'd0;
reg [63:0] storak87 = 64'd0;
reg [63:0] storak88 = 64'd0;
reg [63:0] storak89 = 64'd0;
reg [63:0] storak90 = 64'd0;
reg [63:0] storak91 = 64'd0;
reg [63:0] storak92 = 64'd0;
reg [63:0] storak93 = 64'd0;
reg [63:0] storak94 = 64'd0;
reg [63:0] storak95 = 64'd0;
reg [63:0] storak96 = 64'd0;
reg [63:0] storak97 = 64'd0;
reg [63:0] storak98 = 64'd0;
reg [63:0] storak99 = 64'd0;
reg [63:0] storak100 = 64'd0;
reg [63:0] storak101 = 64'd0;
reg [63:0] storak102 = 64'd0;
reg [63:0] storak103 = 64'd0;
reg [63:0] storak104 = 64'd0;
reg [63:0] storak105 = 64'd0;
reg [63:0] storak106 = 64'd0;
reg [63:0] storak107 = 64'd0;
reg [63:0] storak108 = 64'd0;
reg [63:0] storak109 = 64'd0;
reg [63:0] storak110 = 64'd0;
reg [63:0] storak111 = 64'd0;
reg [63:0] storak112 = 64'd0;
reg [63:0] storak113 = 64'd0;
reg [63:0] storak114 = 64'd0;
reg [63:0] storak115 = 64'd0;
reg [63:0] storak116 = 64'd0;
reg [63:0] storak117 = 64'd0;
reg [63:0] storak118 = 64'd0;
reg [63:0] storak119 = 64'd0;
reg [63:0] storak120 = 64'd0;
reg [63:0] storak121 = 64'd0;
reg [63:0] storak122 = 64'd0;
reg [63:0] storak123 = 64'd0;
reg [63:0] storak124 = 64'd0;
reg [63:0] storak125 = 64'd0;
reg [63:0] storak126 = 64'd0;
reg [63:0] storak127 = 64'd0;
reg [63:0] storav0 = 64'd0;
reg [63:0] storav1 = 64'd0;
reg [63:0] storav2 = 64'd0;
reg [63:0] storav3 = 64'd0;
reg [63:0] storav4 = 64'd0;
reg [63:0] storav5 = 64'd0;
reg [63:0] storav6 = 64'd0;
reg [63:0] storav7 = 64'd0;
reg [63:0] storav8 = 64'd0;
reg [63:0] storav9 = 64'd0;
reg [63:0] storav10 = 64'd0;
reg [63:0] storav11 = 64'd0;
reg [63:0] storav12 = 64'd0;
reg [63:0] storav13 = 64'd0;
reg [63:0] storav14 = 64'd0;
reg [63:0] storav15 = 64'd0;
reg [63:0] storav16 = 64'd0;
reg [63:0] storav17 = 64'd0;
reg [63:0] storav18 = 64'd0;
reg [63:0] storav19 = 64'd0;
reg [63:0] storav20 = 64'd0;
reg [63:0] storav21 = 64'd0;
reg [63:0] storav22 = 64'd0;
reg [63:0] storav23 = 64'd0;
reg [63:0] storav24 = 64'd0;
reg [63:0] storav25 = 64'd0;
reg [63:0] storav26 = 64'd0;
reg [63:0] storav27 = 64'd0;
reg [63:0] storav28 = 64'd0;
reg [63:0] storav29 = 64'd0;
reg [63:0] storav30 = 64'd0;
reg [63:0] storav31 = 64'd0;
reg [63:0] storav32 = 64'd0;
reg [63:0] storav33 = 64'd0;
reg [63:0] storav34 = 64'd0;
reg [63:0] storav35 = 64'd0;
reg [63:0] storav36 = 64'd0;
reg [63:0] storav37 = 64'd0;
reg [63:0] storav38 = 64'd0;
reg [63:0] storav39 = 64'd0;
reg [63:0] storav40 = 64'd0;
reg [63:0] storav41 = 64'd0;
reg [63:0] storav42 = 64'd0;
reg [63:0] storav43 = 64'd0;
reg [63:0] storav44 = 64'd0;
reg [63:0] storav45 = 64'd0;
reg [63:0] storav46 = 64'd0;
reg [63:0] storav47 = 64'd0;
reg [63:0] storav48 = 64'd0;
reg [63:0] storav49 = 64'd0;
reg [63:0] storav50 = 64'd0;
reg [63:0] storav51 = 64'd0;
reg [63:0] storav52 = 64'd0;
reg [63:0] storav53 = 64'd0;
reg [63:0] storav54 = 64'd0;
reg [63:0] storav55 = 64'd0;
reg [63:0] storav56 = 64'd0;
reg [63:0] storav57 = 64'd0;
reg [63:0] storav58 = 64'd0;
reg [63:0] storav59 = 64'd0;
reg [63:0] storav60 = 64'd0;
reg [63:0] storav61 = 64'd0;
reg [63:0] storav62 = 64'd0;
reg [63:0] storav63 = 64'd0;
reg [63:0] storav64 = 64'd0;
reg [63:0] storav65 = 64'd0;
reg [63:0] storav66 = 64'd0;
reg [63:0] storav67 = 64'd0;
reg [63:0] storav68 = 64'd0;
reg [63:0] storav69 = 64'd0;
reg [63:0] storav70 = 64'd0;
reg [63:0] storav71 = 64'd0;
reg [63:0] storav72 = 64'd0;
reg [63:0] storav73 = 64'd0;
reg [63:0] storav74 = 64'd0;
reg [63:0] storav75 = 64'd0;
reg [63:0] storav76 = 64'd0;
reg [63:0] storav77 = 64'd0;
reg [63:0] storav78 = 64'd0;
reg [63:0] storav79 = 64'd0;
reg [63:0] storav80 = 64'd0;
reg [63:0] storav81 = 64'd0;
reg [63:0] storav82 = 64'd0;
reg [63:0] storav83 = 64'd0;
reg [63:0] storav84 = 64'd0;
reg [63:0] storav85 = 64'd0;
reg [63:0] storav86 = 64'd0;
reg [63:0] storav87 = 64'd0;
reg [63:0] storav88 = 64'd0;
reg [63:0] storav89 = 64'd0;
reg [63:0] storav90 = 64'd0;
reg [63:0] storav91 = 64'd0;
reg [63:0] storav92 = 64'd0;
reg [63:0] storav93 = 64'd0;
reg [63:0] storav94 = 64'd0;
reg [63:0] storav95 = 64'd0;
reg [63:0] storav96 = 64'd0;
reg [63:0] storav97 = 64'd0;
reg [63:0] storav98 = 64'd0;
reg [63:0] storav99 = 64'd0;
reg [63:0] storav100 = 64'd0;
reg [63:0] storav101 = 64'd0;
reg [63:0] storav102 = 64'd0;
reg [63:0] storav103 = 64'd0;
reg [63:0] storav104 = 64'd0;
reg [63:0] storav105 = 64'd0;
reg [63:0] storav106 = 64'd0;
reg [63:0] storav107 = 64'd0;
reg [63:0] storav108 = 64'd0;
reg [63:0] storav109 = 64'd0;
reg [63:0] storav110 = 64'd0;
reg [63:0] storav111 = 64'd0;
reg [63:0] storav112 = 64'd0;
reg [63:0] storav113 = 64'd0;
reg [63:0] storav114 = 64'd0;
reg [63:0] storav115 = 64'd0;
reg [63:0] storav116 = 64'd0;
reg [63:0] storav117 = 64'd0;
reg [63:0] storav118 = 64'd0;
reg [63:0] storav119 = 64'd0;
reg [63:0] storav120 = 64'd0;
reg [63:0] storav121 = 64'd0;
reg [63:0] storav122 = 64'd0;
reg [63:0] storav123 = 64'd0;
reg [63:0] storav124 = 64'd0;
reg [63:0] storav125 = 64'd0;
reg [63:0] storav126 = 64'd0;
reg [63:0] storav127 = 64'd0;
reg [63:0] empty_location = 64'd0;
reg [1:0] state = 2'd3;
reg [1:0] next_state;
reg STALL_o_next_value0;
reg STALL_o_next_value_ce0;
reg [63:0] empty_location_t_next_value;
reg empty_location_t_next_value_ce;
reg ACK_o_f_next_value;
reg ACK_o_f_next_value_ce;
reg [63:0] DAT_o_next_value1;
reg DAT_o_next_value_ce1;
reg [63:0] t_next_value0;
reg t_next_value_ce0;
reg [63:0] t_next_value1;
reg t_next_value_ce1;
reg [63:0] f_next_value0;
reg f_next_value_ce0;
reg [63:0] f_next_value1;
reg f_next_value_ce1;
reg [63:0] comb_array_muxed;
reg [63:0] sync_array_muxed0 = 64'd0;
reg [63:0] sync_array_muxed1 = 64'd0;
reg [63:0] sync_array_muxed2 = 64'd0;
reg [63:0] sync_array_muxed3 = 64'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign LA_o = DAT_o;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	next_state <= 2'd0;
	STALL_o_next_value0 <= 1'd0;
	STALL_o_next_value_ce0 <= 1'd0;
	empty_location_t_next_value <= 64'd0;
	empty_location_t_next_value_ce <= 1'd0;
	ACK_o_f_next_value <= 1'd0;
	ACK_o_f_next_value_ce <= 1'd0;
	DAT_o_next_value1 <= 64'd0;
	DAT_o_next_value_ce1 <= 1'd0;
	t_next_value0 <= 64'd0;
	t_next_value_ce0 <= 1'd0;
	t_next_value1 <= 64'd0;
	t_next_value_ce1 <= 1'd0;
	f_next_value0 <= 64'd0;
	f_next_value_ce0 <= 1'd0;
	f_next_value1 <= 64'd0;
	f_next_value_ce1 <= 1'd0;
	next_state <= state;
	case (state)
		1'd0: begin
			STALL_o_next_value0 <= 1'd0;
			STALL_o_next_value_ce0 <= 1'd1;
			if ((((STB_i == 1'd1) & (WE_i == 1'd0)) & (ACK_o == 1'd0))) begin
				next_state <= 1'd1;
			end else begin
				if ((((STB_i == 1'd1) & (WE_i == 1'd1)) & (ACK_o == 1'd0))) begin
					next_state <= 2'd2;
					if ((ADR_i == 64'd0)) begin
						empty_location_t_next_value <= (empty_location + 1'd1);
						empty_location_t_next_value_ce <= 1'd1;
					end
				end else begin
					ACK_o_f_next_value <= 1'd0;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
		end
		1'd1: begin
			if ((ADR_i == 64'd0)) begin
				if ((storak1 == KEY_i)) begin
					DAT_o_next_value1 <= storav1;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak2 == KEY_i)) begin
					DAT_o_next_value1 <= storav2;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak3 == KEY_i)) begin
					DAT_o_next_value1 <= storav3;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak4 == KEY_i)) begin
					DAT_o_next_value1 <= storav4;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak5 == KEY_i)) begin
					DAT_o_next_value1 <= storav5;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak6 == KEY_i)) begin
					DAT_o_next_value1 <= storav6;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak7 == KEY_i)) begin
					DAT_o_next_value1 <= storav7;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak8 == KEY_i)) begin
					DAT_o_next_value1 <= storav8;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak9 == KEY_i)) begin
					DAT_o_next_value1 <= storav9;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak10 == KEY_i)) begin
					DAT_o_next_value1 <= storav10;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak11 == KEY_i)) begin
					DAT_o_next_value1 <= storav11;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak12 == KEY_i)) begin
					DAT_o_next_value1 <= storav12;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak13 == KEY_i)) begin
					DAT_o_next_value1 <= storav13;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak14 == KEY_i)) begin
					DAT_o_next_value1 <= storav14;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak15 == KEY_i)) begin
					DAT_o_next_value1 <= storav15;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak16 == KEY_i)) begin
					DAT_o_next_value1 <= storav16;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak17 == KEY_i)) begin
					DAT_o_next_value1 <= storav17;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak18 == KEY_i)) begin
					DAT_o_next_value1 <= storav18;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak19 == KEY_i)) begin
					DAT_o_next_value1 <= storav19;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak20 == KEY_i)) begin
					DAT_o_next_value1 <= storav20;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak21 == KEY_i)) begin
					DAT_o_next_value1 <= storav21;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak22 == KEY_i)) begin
					DAT_o_next_value1 <= storav22;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak23 == KEY_i)) begin
					DAT_o_next_value1 <= storav23;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak24 == KEY_i)) begin
					DAT_o_next_value1 <= storav24;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak25 == KEY_i)) begin
					DAT_o_next_value1 <= storav25;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak26 == KEY_i)) begin
					DAT_o_next_value1 <= storav26;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak27 == KEY_i)) begin
					DAT_o_next_value1 <= storav27;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak28 == KEY_i)) begin
					DAT_o_next_value1 <= storav28;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak29 == KEY_i)) begin
					DAT_o_next_value1 <= storav29;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak30 == KEY_i)) begin
					DAT_o_next_value1 <= storav30;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak31 == KEY_i)) begin
					DAT_o_next_value1 <= storav31;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak32 == KEY_i)) begin
					DAT_o_next_value1 <= storav32;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak33 == KEY_i)) begin
					DAT_o_next_value1 <= storav33;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak34 == KEY_i)) begin
					DAT_o_next_value1 <= storav34;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak35 == KEY_i)) begin
					DAT_o_next_value1 <= storav35;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak36 == KEY_i)) begin
					DAT_o_next_value1 <= storav36;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak37 == KEY_i)) begin
					DAT_o_next_value1 <= storav37;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak38 == KEY_i)) begin
					DAT_o_next_value1 <= storav38;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak39 == KEY_i)) begin
					DAT_o_next_value1 <= storav39;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak40 == KEY_i)) begin
					DAT_o_next_value1 <= storav40;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak41 == KEY_i)) begin
					DAT_o_next_value1 <= storav41;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak42 == KEY_i)) begin
					DAT_o_next_value1 <= storav42;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak43 == KEY_i)) begin
					DAT_o_next_value1 <= storav43;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak44 == KEY_i)) begin
					DAT_o_next_value1 <= storav44;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak45 == KEY_i)) begin
					DAT_o_next_value1 <= storav45;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak46 == KEY_i)) begin
					DAT_o_next_value1 <= storav46;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak47 == KEY_i)) begin
					DAT_o_next_value1 <= storav47;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak48 == KEY_i)) begin
					DAT_o_next_value1 <= storav48;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak49 == KEY_i)) begin
					DAT_o_next_value1 <= storav49;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak50 == KEY_i)) begin
					DAT_o_next_value1 <= storav50;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak51 == KEY_i)) begin
					DAT_o_next_value1 <= storav51;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak52 == KEY_i)) begin
					DAT_o_next_value1 <= storav52;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak53 == KEY_i)) begin
					DAT_o_next_value1 <= storav53;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak54 == KEY_i)) begin
					DAT_o_next_value1 <= storav54;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak55 == KEY_i)) begin
					DAT_o_next_value1 <= storav55;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak56 == KEY_i)) begin
					DAT_o_next_value1 <= storav56;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak57 == KEY_i)) begin
					DAT_o_next_value1 <= storav57;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak58 == KEY_i)) begin
					DAT_o_next_value1 <= storav58;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak59 == KEY_i)) begin
					DAT_o_next_value1 <= storav59;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak60 == KEY_i)) begin
					DAT_o_next_value1 <= storav60;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak61 == KEY_i)) begin
					DAT_o_next_value1 <= storav61;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak62 == KEY_i)) begin
					DAT_o_next_value1 <= storav62;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak63 == KEY_i)) begin
					DAT_o_next_value1 <= storav63;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak64 == KEY_i)) begin
					DAT_o_next_value1 <= storav64;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak65 == KEY_i)) begin
					DAT_o_next_value1 <= storav65;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak66 == KEY_i)) begin
					DAT_o_next_value1 <= storav66;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak67 == KEY_i)) begin
					DAT_o_next_value1 <= storav67;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak68 == KEY_i)) begin
					DAT_o_next_value1 <= storav68;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak69 == KEY_i)) begin
					DAT_o_next_value1 <= storav69;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak70 == KEY_i)) begin
					DAT_o_next_value1 <= storav70;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak71 == KEY_i)) begin
					DAT_o_next_value1 <= storav71;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak72 == KEY_i)) begin
					DAT_o_next_value1 <= storav72;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak73 == KEY_i)) begin
					DAT_o_next_value1 <= storav73;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak74 == KEY_i)) begin
					DAT_o_next_value1 <= storav74;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak75 == KEY_i)) begin
					DAT_o_next_value1 <= storav75;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak76 == KEY_i)) begin
					DAT_o_next_value1 <= storav76;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak77 == KEY_i)) begin
					DAT_o_next_value1 <= storav77;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak78 == KEY_i)) begin
					DAT_o_next_value1 <= storav78;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak79 == KEY_i)) begin
					DAT_o_next_value1 <= storav79;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak80 == KEY_i)) begin
					DAT_o_next_value1 <= storav80;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak81 == KEY_i)) begin
					DAT_o_next_value1 <= storav81;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak82 == KEY_i)) begin
					DAT_o_next_value1 <= storav82;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak83 == KEY_i)) begin
					DAT_o_next_value1 <= storav83;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak84 == KEY_i)) begin
					DAT_o_next_value1 <= storav84;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak85 == KEY_i)) begin
					DAT_o_next_value1 <= storav85;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak86 == KEY_i)) begin
					DAT_o_next_value1 <= storav86;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak87 == KEY_i)) begin
					DAT_o_next_value1 <= storav87;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak88 == KEY_i)) begin
					DAT_o_next_value1 <= storav88;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak89 == KEY_i)) begin
					DAT_o_next_value1 <= storav89;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak90 == KEY_i)) begin
					DAT_o_next_value1 <= storav90;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak91 == KEY_i)) begin
					DAT_o_next_value1 <= storav91;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak92 == KEY_i)) begin
					DAT_o_next_value1 <= storav92;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak93 == KEY_i)) begin
					DAT_o_next_value1 <= storav93;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak94 == KEY_i)) begin
					DAT_o_next_value1 <= storav94;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak95 == KEY_i)) begin
					DAT_o_next_value1 <= storav95;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak96 == KEY_i)) begin
					DAT_o_next_value1 <= storav96;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak97 == KEY_i)) begin
					DAT_o_next_value1 <= storav97;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak98 == KEY_i)) begin
					DAT_o_next_value1 <= storav98;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak99 == KEY_i)) begin
					DAT_o_next_value1 <= storav99;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak100 == KEY_i)) begin
					DAT_o_next_value1 <= storav100;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak101 == KEY_i)) begin
					DAT_o_next_value1 <= storav101;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak102 == KEY_i)) begin
					DAT_o_next_value1 <= storav102;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak103 == KEY_i)) begin
					DAT_o_next_value1 <= storav103;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak104 == KEY_i)) begin
					DAT_o_next_value1 <= storav104;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak105 == KEY_i)) begin
					DAT_o_next_value1 <= storav105;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak106 == KEY_i)) begin
					DAT_o_next_value1 <= storav106;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak107 == KEY_i)) begin
					DAT_o_next_value1 <= storav107;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak108 == KEY_i)) begin
					DAT_o_next_value1 <= storav108;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak109 == KEY_i)) begin
					DAT_o_next_value1 <= storav109;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak110 == KEY_i)) begin
					DAT_o_next_value1 <= storav110;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak111 == KEY_i)) begin
					DAT_o_next_value1 <= storav111;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak112 == KEY_i)) begin
					DAT_o_next_value1 <= storav112;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak113 == KEY_i)) begin
					DAT_o_next_value1 <= storav113;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak114 == KEY_i)) begin
					DAT_o_next_value1 <= storav114;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak115 == KEY_i)) begin
					DAT_o_next_value1 <= storav115;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak116 == KEY_i)) begin
					DAT_o_next_value1 <= storav116;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak117 == KEY_i)) begin
					DAT_o_next_value1 <= storav117;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak118 == KEY_i)) begin
					DAT_o_next_value1 <= storav118;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak119 == KEY_i)) begin
					DAT_o_next_value1 <= storav119;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak120 == KEY_i)) begin
					DAT_o_next_value1 <= storav120;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak121 == KEY_i)) begin
					DAT_o_next_value1 <= storav121;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak122 == KEY_i)) begin
					DAT_o_next_value1 <= storav122;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak123 == KEY_i)) begin
					DAT_o_next_value1 <= storav123;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak124 == KEY_i)) begin
					DAT_o_next_value1 <= storav124;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak125 == KEY_i)) begin
					DAT_o_next_value1 <= storav125;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak126 == KEY_i)) begin
					DAT_o_next_value1 <= storav126;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i == 64'd0)) begin
				if ((storak127 == KEY_i)) begin
					DAT_o_next_value1 <= storav127;
					DAT_o_next_value_ce1 <= 1'd1;
					ACK_o_f_next_value <= 1'd1;
					ACK_o_f_next_value_ce <= 1'd1;
					next_state <= 1'd0;
				end
			end
			if ((ADR_i != 64'd0)) begin
				DAT_o_next_value1 <= comb_array_muxed;
				DAT_o_next_value_ce1 <= 1'd1;
				ACK_o_f_next_value <= 1'd1;
				ACK_o_f_next_value_ce <= 1'd1;
				next_state <= 1'd0;
			end
			if ((sys_rst == 1'd1)) begin
				next_state <= 2'd3;
			end
		end
		2'd2: begin
			if ((ADR_i == 64'd0)) begin
				t_next_value0 <= DAT_i;
				t_next_value_ce0 <= 1'd1;
				t_next_value1 <= KEY_i;
				t_next_value_ce1 <= 1'd1;
				DAT_o_next_value1 <= empty_location;
				DAT_o_next_value_ce1 <= 1'd1;
			end else begin
				f_next_value0 <= DAT_i;
				f_next_value_ce0 <= 1'd1;
				f_next_value1 <= KEY_i;
				f_next_value_ce1 <= 1'd1;
				DAT_o_next_value1 <= ADR_i;
				DAT_o_next_value_ce1 <= 1'd1;
			end
			ACK_o_f_next_value <= 1'd1;
			ACK_o_f_next_value_ce <= 1'd1;
			next_state <= 1'd0;
			if ((sys_rst == 1'd1)) begin
				next_state <= 2'd3;
			end else begin
				next_state <= 1'd0;
			end
		end
		default: begin
			next_state <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	comb_array_muxed <= 64'd0;
	case (ADR_i)
		1'd0: begin
			comb_array_muxed <= storav0;
		end
		1'd1: begin
			comb_array_muxed <= storav1;
		end
		2'd2: begin
			comb_array_muxed <= storav2;
		end
		2'd3: begin
			comb_array_muxed <= storav3;
		end
		3'd4: begin
			comb_array_muxed <= storav4;
		end
		3'd5: begin
			comb_array_muxed <= storav5;
		end
		3'd6: begin
			comb_array_muxed <= storav6;
		end
		3'd7: begin
			comb_array_muxed <= storav7;
		end
		4'd8: begin
			comb_array_muxed <= storav8;
		end
		4'd9: begin
			comb_array_muxed <= storav9;
		end
		4'd10: begin
			comb_array_muxed <= storav10;
		end
		4'd11: begin
			comb_array_muxed <= storav11;
		end
		4'd12: begin
			comb_array_muxed <= storav12;
		end
		4'd13: begin
			comb_array_muxed <= storav13;
		end
		4'd14: begin
			comb_array_muxed <= storav14;
		end
		4'd15: begin
			comb_array_muxed <= storav15;
		end
		5'd16: begin
			comb_array_muxed <= storav16;
		end
		5'd17: begin
			comb_array_muxed <= storav17;
		end
		5'd18: begin
			comb_array_muxed <= storav18;
		end
		5'd19: begin
			comb_array_muxed <= storav19;
		end
		5'd20: begin
			comb_array_muxed <= storav20;
		end
		5'd21: begin
			comb_array_muxed <= storav21;
		end
		5'd22: begin
			comb_array_muxed <= storav22;
		end
		5'd23: begin
			comb_array_muxed <= storav23;
		end
		5'd24: begin
			comb_array_muxed <= storav24;
		end
		5'd25: begin
			comb_array_muxed <= storav25;
		end
		5'd26: begin
			comb_array_muxed <= storav26;
		end
		5'd27: begin
			comb_array_muxed <= storav27;
		end
		5'd28: begin
			comb_array_muxed <= storav28;
		end
		5'd29: begin
			comb_array_muxed <= storav29;
		end
		5'd30: begin
			comb_array_muxed <= storav30;
		end
		5'd31: begin
			comb_array_muxed <= storav31;
		end
		6'd32: begin
			comb_array_muxed <= storav32;
		end
		6'd33: begin
			comb_array_muxed <= storav33;
		end
		6'd34: begin
			comb_array_muxed <= storav34;
		end
		6'd35: begin
			comb_array_muxed <= storav35;
		end
		6'd36: begin
			comb_array_muxed <= storav36;
		end
		6'd37: begin
			comb_array_muxed <= storav37;
		end
		6'd38: begin
			comb_array_muxed <= storav38;
		end
		6'd39: begin
			comb_array_muxed <= storav39;
		end
		6'd40: begin
			comb_array_muxed <= storav40;
		end
		6'd41: begin
			comb_array_muxed <= storav41;
		end
		6'd42: begin
			comb_array_muxed <= storav42;
		end
		6'd43: begin
			comb_array_muxed <= storav43;
		end
		6'd44: begin
			comb_array_muxed <= storav44;
		end
		6'd45: begin
			comb_array_muxed <= storav45;
		end
		6'd46: begin
			comb_array_muxed <= storav46;
		end
		6'd47: begin
			comb_array_muxed <= storav47;
		end
		6'd48: begin
			comb_array_muxed <= storav48;
		end
		6'd49: begin
			comb_array_muxed <= storav49;
		end
		6'd50: begin
			comb_array_muxed <= storav50;
		end
		6'd51: begin
			comb_array_muxed <= storav51;
		end
		6'd52: begin
			comb_array_muxed <= storav52;
		end
		6'd53: begin
			comb_array_muxed <= storav53;
		end
		6'd54: begin
			comb_array_muxed <= storav54;
		end
		6'd55: begin
			comb_array_muxed <= storav55;
		end
		6'd56: begin
			comb_array_muxed <= storav56;
		end
		6'd57: begin
			comb_array_muxed <= storav57;
		end
		6'd58: begin
			comb_array_muxed <= storav58;
		end
		6'd59: begin
			comb_array_muxed <= storav59;
		end
		6'd60: begin
			comb_array_muxed <= storav60;
		end
		6'd61: begin
			comb_array_muxed <= storav61;
		end
		6'd62: begin
			comb_array_muxed <= storav62;
		end
		6'd63: begin
			comb_array_muxed <= storav63;
		end
		7'd64: begin
			comb_array_muxed <= storav64;
		end
		7'd65: begin
			comb_array_muxed <= storav65;
		end
		7'd66: begin
			comb_array_muxed <= storav66;
		end
		7'd67: begin
			comb_array_muxed <= storav67;
		end
		7'd68: begin
			comb_array_muxed <= storav68;
		end
		7'd69: begin
			comb_array_muxed <= storav69;
		end
		7'd70: begin
			comb_array_muxed <= storav70;
		end
		7'd71: begin
			comb_array_muxed <= storav71;
		end
		7'd72: begin
			comb_array_muxed <= storav72;
		end
		7'd73: begin
			comb_array_muxed <= storav73;
		end
		7'd74: begin
			comb_array_muxed <= storav74;
		end
		7'd75: begin
			comb_array_muxed <= storav75;
		end
		7'd76: begin
			comb_array_muxed <= storav76;
		end
		7'd77: begin
			comb_array_muxed <= storav77;
		end
		7'd78: begin
			comb_array_muxed <= storav78;
		end
		7'd79: begin
			comb_array_muxed <= storav79;
		end
		7'd80: begin
			comb_array_muxed <= storav80;
		end
		7'd81: begin
			comb_array_muxed <= storav81;
		end
		7'd82: begin
			comb_array_muxed <= storav82;
		end
		7'd83: begin
			comb_array_muxed <= storav83;
		end
		7'd84: begin
			comb_array_muxed <= storav84;
		end
		7'd85: begin
			comb_array_muxed <= storav85;
		end
		7'd86: begin
			comb_array_muxed <= storav86;
		end
		7'd87: begin
			comb_array_muxed <= storav87;
		end
		7'd88: begin
			comb_array_muxed <= storav88;
		end
		7'd89: begin
			comb_array_muxed <= storav89;
		end
		7'd90: begin
			comb_array_muxed <= storav90;
		end
		7'd91: begin
			comb_array_muxed <= storav91;
		end
		7'd92: begin
			comb_array_muxed <= storav92;
		end
		7'd93: begin
			comb_array_muxed <= storav93;
		end
		7'd94: begin
			comb_array_muxed <= storav94;
		end
		7'd95: begin
			comb_array_muxed <= storav95;
		end
		7'd96: begin
			comb_array_muxed <= storav96;
		end
		7'd97: begin
			comb_array_muxed <= storav97;
		end
		7'd98: begin
			comb_array_muxed <= storav98;
		end
		7'd99: begin
			comb_array_muxed <= storav99;
		end
		7'd100: begin
			comb_array_muxed <= storav100;
		end
		7'd101: begin
			comb_array_muxed <= storav101;
		end
		7'd102: begin
			comb_array_muxed <= storav102;
		end
		7'd103: begin
			comb_array_muxed <= storav103;
		end
		7'd104: begin
			comb_array_muxed <= storav104;
		end
		7'd105: begin
			comb_array_muxed <= storav105;
		end
		7'd106: begin
			comb_array_muxed <= storav106;
		end
		7'd107: begin
			comb_array_muxed <= storav107;
		end
		7'd108: begin
			comb_array_muxed <= storav108;
		end
		7'd109: begin
			comb_array_muxed <= storav109;
		end
		7'd110: begin
			comb_array_muxed <= storav110;
		end
		7'd111: begin
			comb_array_muxed <= storav111;
		end
		7'd112: begin
			comb_array_muxed <= storav112;
		end
		7'd113: begin
			comb_array_muxed <= storav113;
		end
		7'd114: begin
			comb_array_muxed <= storav114;
		end
		7'd115: begin
			comb_array_muxed <= storav115;
		end
		7'd116: begin
			comb_array_muxed <= storav116;
		end
		7'd117: begin
			comb_array_muxed <= storav117;
		end
		7'd118: begin
			comb_array_muxed <= storav118;
		end
		7'd119: begin
			comb_array_muxed <= storav119;
		end
		7'd120: begin
			comb_array_muxed <= storav120;
		end
		7'd121: begin
			comb_array_muxed <= storav121;
		end
		7'd122: begin
			comb_array_muxed <= storav122;
		end
		7'd123: begin
			comb_array_muxed <= storav123;
		end
		7'd124: begin
			comb_array_muxed <= storav124;
		end
		7'd125: begin
			comb_array_muxed <= storav125;
		end
		7'd126: begin
			comb_array_muxed <= storav126;
		end
		default: begin
			comb_array_muxed <= storav127;
		end
	endcase
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

always @(posedge sys_clk) begin
	state <= next_state;
	if (STALL_o_next_value_ce0) begin
		STALL_o <= STALL_o_next_value0;
	end
	if (empty_location_t_next_value_ce) begin
		empty_location <= empty_location_t_next_value;
	end
	if (ACK_o_f_next_value_ce) begin
		ACK_o <= ACK_o_f_next_value;
	end
	if (DAT_o_next_value_ce1) begin
		DAT_o <= DAT_o_next_value1;
	end
	if (t_next_value_ce0) begin
		sync_array_muxed0 = t_next_value0;
		case (empty_location)
			1'd0: begin
				storav0 <= sync_array_muxed0;
			end
			1'd1: begin
				storav1 <= sync_array_muxed0;
			end
			2'd2: begin
				storav2 <= sync_array_muxed0;
			end
			2'd3: begin
				storav3 <= sync_array_muxed0;
			end
			3'd4: begin
				storav4 <= sync_array_muxed0;
			end
			3'd5: begin
				storav5 <= sync_array_muxed0;
			end
			3'd6: begin
				storav6 <= sync_array_muxed0;
			end
			3'd7: begin
				storav7 <= sync_array_muxed0;
			end
			4'd8: begin
				storav8 <= sync_array_muxed0;
			end
			4'd9: begin
				storav9 <= sync_array_muxed0;
			end
			4'd10: begin
				storav10 <= sync_array_muxed0;
			end
			4'd11: begin
				storav11 <= sync_array_muxed0;
			end
			4'd12: begin
				storav12 <= sync_array_muxed0;
			end
			4'd13: begin
				storav13 <= sync_array_muxed0;
			end
			4'd14: begin
				storav14 <= sync_array_muxed0;
			end
			4'd15: begin
				storav15 <= sync_array_muxed0;
			end
			5'd16: begin
				storav16 <= sync_array_muxed0;
			end
			5'd17: begin
				storav17 <= sync_array_muxed0;
			end
			5'd18: begin
				storav18 <= sync_array_muxed0;
			end
			5'd19: begin
				storav19 <= sync_array_muxed0;
			end
			5'd20: begin
				storav20 <= sync_array_muxed0;
			end
			5'd21: begin
				storav21 <= sync_array_muxed0;
			end
			5'd22: begin
				storav22 <= sync_array_muxed0;
			end
			5'd23: begin
				storav23 <= sync_array_muxed0;
			end
			5'd24: begin
				storav24 <= sync_array_muxed0;
			end
			5'd25: begin
				storav25 <= sync_array_muxed0;
			end
			5'd26: begin
				storav26 <= sync_array_muxed0;
			end
			5'd27: begin
				storav27 <= sync_array_muxed0;
			end
			5'd28: begin
				storav28 <= sync_array_muxed0;
			end
			5'd29: begin
				storav29 <= sync_array_muxed0;
			end
			5'd30: begin
				storav30 <= sync_array_muxed0;
			end
			5'd31: begin
				storav31 <= sync_array_muxed0;
			end
			6'd32: begin
				storav32 <= sync_array_muxed0;
			end
			6'd33: begin
				storav33 <= sync_array_muxed0;
			end
			6'd34: begin
				storav34 <= sync_array_muxed0;
			end
			6'd35: begin
				storav35 <= sync_array_muxed0;
			end
			6'd36: begin
				storav36 <= sync_array_muxed0;
			end
			6'd37: begin
				storav37 <= sync_array_muxed0;
			end
			6'd38: begin
				storav38 <= sync_array_muxed0;
			end
			6'd39: begin
				storav39 <= sync_array_muxed0;
			end
			6'd40: begin
				storav40 <= sync_array_muxed0;
			end
			6'd41: begin
				storav41 <= sync_array_muxed0;
			end
			6'd42: begin
				storav42 <= sync_array_muxed0;
			end
			6'd43: begin
				storav43 <= sync_array_muxed0;
			end
			6'd44: begin
				storav44 <= sync_array_muxed0;
			end
			6'd45: begin
				storav45 <= sync_array_muxed0;
			end
			6'd46: begin
				storav46 <= sync_array_muxed0;
			end
			6'd47: begin
				storav47 <= sync_array_muxed0;
			end
			6'd48: begin
				storav48 <= sync_array_muxed0;
			end
			6'd49: begin
				storav49 <= sync_array_muxed0;
			end
			6'd50: begin
				storav50 <= sync_array_muxed0;
			end
			6'd51: begin
				storav51 <= sync_array_muxed0;
			end
			6'd52: begin
				storav52 <= sync_array_muxed0;
			end
			6'd53: begin
				storav53 <= sync_array_muxed0;
			end
			6'd54: begin
				storav54 <= sync_array_muxed0;
			end
			6'd55: begin
				storav55 <= sync_array_muxed0;
			end
			6'd56: begin
				storav56 <= sync_array_muxed0;
			end
			6'd57: begin
				storav57 <= sync_array_muxed0;
			end
			6'd58: begin
				storav58 <= sync_array_muxed0;
			end
			6'd59: begin
				storav59 <= sync_array_muxed0;
			end
			6'd60: begin
				storav60 <= sync_array_muxed0;
			end
			6'd61: begin
				storav61 <= sync_array_muxed0;
			end
			6'd62: begin
				storav62 <= sync_array_muxed0;
			end
			6'd63: begin
				storav63 <= sync_array_muxed0;
			end
			7'd64: begin
				storav64 <= sync_array_muxed0;
			end
			7'd65: begin
				storav65 <= sync_array_muxed0;
			end
			7'd66: begin
				storav66 <= sync_array_muxed0;
			end
			7'd67: begin
				storav67 <= sync_array_muxed0;
			end
			7'd68: begin
				storav68 <= sync_array_muxed0;
			end
			7'd69: begin
				storav69 <= sync_array_muxed0;
			end
			7'd70: begin
				storav70 <= sync_array_muxed0;
			end
			7'd71: begin
				storav71 <= sync_array_muxed0;
			end
			7'd72: begin
				storav72 <= sync_array_muxed0;
			end
			7'd73: begin
				storav73 <= sync_array_muxed0;
			end
			7'd74: begin
				storav74 <= sync_array_muxed0;
			end
			7'd75: begin
				storav75 <= sync_array_muxed0;
			end
			7'd76: begin
				storav76 <= sync_array_muxed0;
			end
			7'd77: begin
				storav77 <= sync_array_muxed0;
			end
			7'd78: begin
				storav78 <= sync_array_muxed0;
			end
			7'd79: begin
				storav79 <= sync_array_muxed0;
			end
			7'd80: begin
				storav80 <= sync_array_muxed0;
			end
			7'd81: begin
				storav81 <= sync_array_muxed0;
			end
			7'd82: begin
				storav82 <= sync_array_muxed0;
			end
			7'd83: begin
				storav83 <= sync_array_muxed0;
			end
			7'd84: begin
				storav84 <= sync_array_muxed0;
			end
			7'd85: begin
				storav85 <= sync_array_muxed0;
			end
			7'd86: begin
				storav86 <= sync_array_muxed0;
			end
			7'd87: begin
				storav87 <= sync_array_muxed0;
			end
			7'd88: begin
				storav88 <= sync_array_muxed0;
			end
			7'd89: begin
				storav89 <= sync_array_muxed0;
			end
			7'd90: begin
				storav90 <= sync_array_muxed0;
			end
			7'd91: begin
				storav91 <= sync_array_muxed0;
			end
			7'd92: begin
				storav92 <= sync_array_muxed0;
			end
			7'd93: begin
				storav93 <= sync_array_muxed0;
			end
			7'd94: begin
				storav94 <= sync_array_muxed0;
			end
			7'd95: begin
				storav95 <= sync_array_muxed0;
			end
			7'd96: begin
				storav96 <= sync_array_muxed0;
			end
			7'd97: begin
				storav97 <= sync_array_muxed0;
			end
			7'd98: begin
				storav98 <= sync_array_muxed0;
			end
			7'd99: begin
				storav99 <= sync_array_muxed0;
			end
			7'd100: begin
				storav100 <= sync_array_muxed0;
			end
			7'd101: begin
				storav101 <= sync_array_muxed0;
			end
			7'd102: begin
				storav102 <= sync_array_muxed0;
			end
			7'd103: begin
				storav103 <= sync_array_muxed0;
			end
			7'd104: begin
				storav104 <= sync_array_muxed0;
			end
			7'd105: begin
				storav105 <= sync_array_muxed0;
			end
			7'd106: begin
				storav106 <= sync_array_muxed0;
			end
			7'd107: begin
				storav107 <= sync_array_muxed0;
			end
			7'd108: begin
				storav108 <= sync_array_muxed0;
			end
			7'd109: begin
				storav109 <= sync_array_muxed0;
			end
			7'd110: begin
				storav110 <= sync_array_muxed0;
			end
			7'd111: begin
				storav111 <= sync_array_muxed0;
			end
			7'd112: begin
				storav112 <= sync_array_muxed0;
			end
			7'd113: begin
				storav113 <= sync_array_muxed0;
			end
			7'd114: begin
				storav114 <= sync_array_muxed0;
			end
			7'd115: begin
				storav115 <= sync_array_muxed0;
			end
			7'd116: begin
				storav116 <= sync_array_muxed0;
			end
			7'd117: begin
				storav117 <= sync_array_muxed0;
			end
			7'd118: begin
				storav118 <= sync_array_muxed0;
			end
			7'd119: begin
				storav119 <= sync_array_muxed0;
			end
			7'd120: begin
				storav120 <= sync_array_muxed0;
			end
			7'd121: begin
				storav121 <= sync_array_muxed0;
			end
			7'd122: begin
				storav122 <= sync_array_muxed0;
			end
			7'd123: begin
				storav123 <= sync_array_muxed0;
			end
			7'd124: begin
				storav124 <= sync_array_muxed0;
			end
			7'd125: begin
				storav125 <= sync_array_muxed0;
			end
			7'd126: begin
				storav126 <= sync_array_muxed0;
			end
			default: begin
				storav127 <= sync_array_muxed0;
			end
		endcase
	end
	if (t_next_value_ce1) begin
		sync_array_muxed1 = t_next_value1;
		case (empty_location)
			1'd0: begin
				storak0 <= sync_array_muxed1;
			end
			1'd1: begin
				storak1 <= sync_array_muxed1;
			end
			2'd2: begin
				storak2 <= sync_array_muxed1;
			end
			2'd3: begin
				storak3 <= sync_array_muxed1;
			end
			3'd4: begin
				storak4 <= sync_array_muxed1;
			end
			3'd5: begin
				storak5 <= sync_array_muxed1;
			end
			3'd6: begin
				storak6 <= sync_array_muxed1;
			end
			3'd7: begin
				storak7 <= sync_array_muxed1;
			end
			4'd8: begin
				storak8 <= sync_array_muxed1;
			end
			4'd9: begin
				storak9 <= sync_array_muxed1;
			end
			4'd10: begin
				storak10 <= sync_array_muxed1;
			end
			4'd11: begin
				storak11 <= sync_array_muxed1;
			end
			4'd12: begin
				storak12 <= sync_array_muxed1;
			end
			4'd13: begin
				storak13 <= sync_array_muxed1;
			end
			4'd14: begin
				storak14 <= sync_array_muxed1;
			end
			4'd15: begin
				storak15 <= sync_array_muxed1;
			end
			5'd16: begin
				storak16 <= sync_array_muxed1;
			end
			5'd17: begin
				storak17 <= sync_array_muxed1;
			end
			5'd18: begin
				storak18 <= sync_array_muxed1;
			end
			5'd19: begin
				storak19 <= sync_array_muxed1;
			end
			5'd20: begin
				storak20 <= sync_array_muxed1;
			end
			5'd21: begin
				storak21 <= sync_array_muxed1;
			end
			5'd22: begin
				storak22 <= sync_array_muxed1;
			end
			5'd23: begin
				storak23 <= sync_array_muxed1;
			end
			5'd24: begin
				storak24 <= sync_array_muxed1;
			end
			5'd25: begin
				storak25 <= sync_array_muxed1;
			end
			5'd26: begin
				storak26 <= sync_array_muxed1;
			end
			5'd27: begin
				storak27 <= sync_array_muxed1;
			end
			5'd28: begin
				storak28 <= sync_array_muxed1;
			end
			5'd29: begin
				storak29 <= sync_array_muxed1;
			end
			5'd30: begin
				storak30 <= sync_array_muxed1;
			end
			5'd31: begin
				storak31 <= sync_array_muxed1;
			end
			6'd32: begin
				storak32 <= sync_array_muxed1;
			end
			6'd33: begin
				storak33 <= sync_array_muxed1;
			end
			6'd34: begin
				storak34 <= sync_array_muxed1;
			end
			6'd35: begin
				storak35 <= sync_array_muxed1;
			end
			6'd36: begin
				storak36 <= sync_array_muxed1;
			end
			6'd37: begin
				storak37 <= sync_array_muxed1;
			end
			6'd38: begin
				storak38 <= sync_array_muxed1;
			end
			6'd39: begin
				storak39 <= sync_array_muxed1;
			end
			6'd40: begin
				storak40 <= sync_array_muxed1;
			end
			6'd41: begin
				storak41 <= sync_array_muxed1;
			end
			6'd42: begin
				storak42 <= sync_array_muxed1;
			end
			6'd43: begin
				storak43 <= sync_array_muxed1;
			end
			6'd44: begin
				storak44 <= sync_array_muxed1;
			end
			6'd45: begin
				storak45 <= sync_array_muxed1;
			end
			6'd46: begin
				storak46 <= sync_array_muxed1;
			end
			6'd47: begin
				storak47 <= sync_array_muxed1;
			end
			6'd48: begin
				storak48 <= sync_array_muxed1;
			end
			6'd49: begin
				storak49 <= sync_array_muxed1;
			end
			6'd50: begin
				storak50 <= sync_array_muxed1;
			end
			6'd51: begin
				storak51 <= sync_array_muxed1;
			end
			6'd52: begin
				storak52 <= sync_array_muxed1;
			end
			6'd53: begin
				storak53 <= sync_array_muxed1;
			end
			6'd54: begin
				storak54 <= sync_array_muxed1;
			end
			6'd55: begin
				storak55 <= sync_array_muxed1;
			end
			6'd56: begin
				storak56 <= sync_array_muxed1;
			end
			6'd57: begin
				storak57 <= sync_array_muxed1;
			end
			6'd58: begin
				storak58 <= sync_array_muxed1;
			end
			6'd59: begin
				storak59 <= sync_array_muxed1;
			end
			6'd60: begin
				storak60 <= sync_array_muxed1;
			end
			6'd61: begin
				storak61 <= sync_array_muxed1;
			end
			6'd62: begin
				storak62 <= sync_array_muxed1;
			end
			6'd63: begin
				storak63 <= sync_array_muxed1;
			end
			7'd64: begin
				storak64 <= sync_array_muxed1;
			end
			7'd65: begin
				storak65 <= sync_array_muxed1;
			end
			7'd66: begin
				storak66 <= sync_array_muxed1;
			end
			7'd67: begin
				storak67 <= sync_array_muxed1;
			end
			7'd68: begin
				storak68 <= sync_array_muxed1;
			end
			7'd69: begin
				storak69 <= sync_array_muxed1;
			end
			7'd70: begin
				storak70 <= sync_array_muxed1;
			end
			7'd71: begin
				storak71 <= sync_array_muxed1;
			end
			7'd72: begin
				storak72 <= sync_array_muxed1;
			end
			7'd73: begin
				storak73 <= sync_array_muxed1;
			end
			7'd74: begin
				storak74 <= sync_array_muxed1;
			end
			7'd75: begin
				storak75 <= sync_array_muxed1;
			end
			7'd76: begin
				storak76 <= sync_array_muxed1;
			end
			7'd77: begin
				storak77 <= sync_array_muxed1;
			end
			7'd78: begin
				storak78 <= sync_array_muxed1;
			end
			7'd79: begin
				storak79 <= sync_array_muxed1;
			end
			7'd80: begin
				storak80 <= sync_array_muxed1;
			end
			7'd81: begin
				storak81 <= sync_array_muxed1;
			end
			7'd82: begin
				storak82 <= sync_array_muxed1;
			end
			7'd83: begin
				storak83 <= sync_array_muxed1;
			end
			7'd84: begin
				storak84 <= sync_array_muxed1;
			end
			7'd85: begin
				storak85 <= sync_array_muxed1;
			end
			7'd86: begin
				storak86 <= sync_array_muxed1;
			end
			7'd87: begin
				storak87 <= sync_array_muxed1;
			end
			7'd88: begin
				storak88 <= sync_array_muxed1;
			end
			7'd89: begin
				storak89 <= sync_array_muxed1;
			end
			7'd90: begin
				storak90 <= sync_array_muxed1;
			end
			7'd91: begin
				storak91 <= sync_array_muxed1;
			end
			7'd92: begin
				storak92 <= sync_array_muxed1;
			end
			7'd93: begin
				storak93 <= sync_array_muxed1;
			end
			7'd94: begin
				storak94 <= sync_array_muxed1;
			end
			7'd95: begin
				storak95 <= sync_array_muxed1;
			end
			7'd96: begin
				storak96 <= sync_array_muxed1;
			end
			7'd97: begin
				storak97 <= sync_array_muxed1;
			end
			7'd98: begin
				storak98 <= sync_array_muxed1;
			end
			7'd99: begin
				storak99 <= sync_array_muxed1;
			end
			7'd100: begin
				storak100 <= sync_array_muxed1;
			end
			7'd101: begin
				storak101 <= sync_array_muxed1;
			end
			7'd102: begin
				storak102 <= sync_array_muxed1;
			end
			7'd103: begin
				storak103 <= sync_array_muxed1;
			end
			7'd104: begin
				storak104 <= sync_array_muxed1;
			end
			7'd105: begin
				storak105 <= sync_array_muxed1;
			end
			7'd106: begin
				storak106 <= sync_array_muxed1;
			end
			7'd107: begin
				storak107 <= sync_array_muxed1;
			end
			7'd108: begin
				storak108 <= sync_array_muxed1;
			end
			7'd109: begin
				storak109 <= sync_array_muxed1;
			end
			7'd110: begin
				storak110 <= sync_array_muxed1;
			end
			7'd111: begin
				storak111 <= sync_array_muxed1;
			end
			7'd112: begin
				storak112 <= sync_array_muxed1;
			end
			7'd113: begin
				storak113 <= sync_array_muxed1;
			end
			7'd114: begin
				storak114 <= sync_array_muxed1;
			end
			7'd115: begin
				storak115 <= sync_array_muxed1;
			end
			7'd116: begin
				storak116 <= sync_array_muxed1;
			end
			7'd117: begin
				storak117 <= sync_array_muxed1;
			end
			7'd118: begin
				storak118 <= sync_array_muxed1;
			end
			7'd119: begin
				storak119 <= sync_array_muxed1;
			end
			7'd120: begin
				storak120 <= sync_array_muxed1;
			end
			7'd121: begin
				storak121 <= sync_array_muxed1;
			end
			7'd122: begin
				storak122 <= sync_array_muxed1;
			end
			7'd123: begin
				storak123 <= sync_array_muxed1;
			end
			7'd124: begin
				storak124 <= sync_array_muxed1;
			end
			7'd125: begin
				storak125 <= sync_array_muxed1;
			end
			7'd126: begin
				storak126 <= sync_array_muxed1;
			end
			default: begin
				storak127 <= sync_array_muxed1;
			end
		endcase
	end
	if (f_next_value_ce0) begin
		sync_array_muxed2 = f_next_value0;
		case (ADR_i)
			1'd0: begin
				storav0 <= sync_array_muxed2;
			end
			1'd1: begin
				storav1 <= sync_array_muxed2;
			end
			2'd2: begin
				storav2 <= sync_array_muxed2;
			end
			2'd3: begin
				storav3 <= sync_array_muxed2;
			end
			3'd4: begin
				storav4 <= sync_array_muxed2;
			end
			3'd5: begin
				storav5 <= sync_array_muxed2;
			end
			3'd6: begin
				storav6 <= sync_array_muxed2;
			end
			3'd7: begin
				storav7 <= sync_array_muxed2;
			end
			4'd8: begin
				storav8 <= sync_array_muxed2;
			end
			4'd9: begin
				storav9 <= sync_array_muxed2;
			end
			4'd10: begin
				storav10 <= sync_array_muxed2;
			end
			4'd11: begin
				storav11 <= sync_array_muxed2;
			end
			4'd12: begin
				storav12 <= sync_array_muxed2;
			end
			4'd13: begin
				storav13 <= sync_array_muxed2;
			end
			4'd14: begin
				storav14 <= sync_array_muxed2;
			end
			4'd15: begin
				storav15 <= sync_array_muxed2;
			end
			5'd16: begin
				storav16 <= sync_array_muxed2;
			end
			5'd17: begin
				storav17 <= sync_array_muxed2;
			end
			5'd18: begin
				storav18 <= sync_array_muxed2;
			end
			5'd19: begin
				storav19 <= sync_array_muxed2;
			end
			5'd20: begin
				storav20 <= sync_array_muxed2;
			end
			5'd21: begin
				storav21 <= sync_array_muxed2;
			end
			5'd22: begin
				storav22 <= sync_array_muxed2;
			end
			5'd23: begin
				storav23 <= sync_array_muxed2;
			end
			5'd24: begin
				storav24 <= sync_array_muxed2;
			end
			5'd25: begin
				storav25 <= sync_array_muxed2;
			end
			5'd26: begin
				storav26 <= sync_array_muxed2;
			end
			5'd27: begin
				storav27 <= sync_array_muxed2;
			end
			5'd28: begin
				storav28 <= sync_array_muxed2;
			end
			5'd29: begin
				storav29 <= sync_array_muxed2;
			end
			5'd30: begin
				storav30 <= sync_array_muxed2;
			end
			5'd31: begin
				storav31 <= sync_array_muxed2;
			end
			6'd32: begin
				storav32 <= sync_array_muxed2;
			end
			6'd33: begin
				storav33 <= sync_array_muxed2;
			end
			6'd34: begin
				storav34 <= sync_array_muxed2;
			end
			6'd35: begin
				storav35 <= sync_array_muxed2;
			end
			6'd36: begin
				storav36 <= sync_array_muxed2;
			end
			6'd37: begin
				storav37 <= sync_array_muxed2;
			end
			6'd38: begin
				storav38 <= sync_array_muxed2;
			end
			6'd39: begin
				storav39 <= sync_array_muxed2;
			end
			6'd40: begin
				storav40 <= sync_array_muxed2;
			end
			6'd41: begin
				storav41 <= sync_array_muxed2;
			end
			6'd42: begin
				storav42 <= sync_array_muxed2;
			end
			6'd43: begin
				storav43 <= sync_array_muxed2;
			end
			6'd44: begin
				storav44 <= sync_array_muxed2;
			end
			6'd45: begin
				storav45 <= sync_array_muxed2;
			end
			6'd46: begin
				storav46 <= sync_array_muxed2;
			end
			6'd47: begin
				storav47 <= sync_array_muxed2;
			end
			6'd48: begin
				storav48 <= sync_array_muxed2;
			end
			6'd49: begin
				storav49 <= sync_array_muxed2;
			end
			6'd50: begin
				storav50 <= sync_array_muxed2;
			end
			6'd51: begin
				storav51 <= sync_array_muxed2;
			end
			6'd52: begin
				storav52 <= sync_array_muxed2;
			end
			6'd53: begin
				storav53 <= sync_array_muxed2;
			end
			6'd54: begin
				storav54 <= sync_array_muxed2;
			end
			6'd55: begin
				storav55 <= sync_array_muxed2;
			end
			6'd56: begin
				storav56 <= sync_array_muxed2;
			end
			6'd57: begin
				storav57 <= sync_array_muxed2;
			end
			6'd58: begin
				storav58 <= sync_array_muxed2;
			end
			6'd59: begin
				storav59 <= sync_array_muxed2;
			end
			6'd60: begin
				storav60 <= sync_array_muxed2;
			end
			6'd61: begin
				storav61 <= sync_array_muxed2;
			end
			6'd62: begin
				storav62 <= sync_array_muxed2;
			end
			6'd63: begin
				storav63 <= sync_array_muxed2;
			end
			7'd64: begin
				storav64 <= sync_array_muxed2;
			end
			7'd65: begin
				storav65 <= sync_array_muxed2;
			end
			7'd66: begin
				storav66 <= sync_array_muxed2;
			end
			7'd67: begin
				storav67 <= sync_array_muxed2;
			end
			7'd68: begin
				storav68 <= sync_array_muxed2;
			end
			7'd69: begin
				storav69 <= sync_array_muxed2;
			end
			7'd70: begin
				storav70 <= sync_array_muxed2;
			end
			7'd71: begin
				storav71 <= sync_array_muxed2;
			end
			7'd72: begin
				storav72 <= sync_array_muxed2;
			end
			7'd73: begin
				storav73 <= sync_array_muxed2;
			end
			7'd74: begin
				storav74 <= sync_array_muxed2;
			end
			7'd75: begin
				storav75 <= sync_array_muxed2;
			end
			7'd76: begin
				storav76 <= sync_array_muxed2;
			end
			7'd77: begin
				storav77 <= sync_array_muxed2;
			end
			7'd78: begin
				storav78 <= sync_array_muxed2;
			end
			7'd79: begin
				storav79 <= sync_array_muxed2;
			end
			7'd80: begin
				storav80 <= sync_array_muxed2;
			end
			7'd81: begin
				storav81 <= sync_array_muxed2;
			end
			7'd82: begin
				storav82 <= sync_array_muxed2;
			end
			7'd83: begin
				storav83 <= sync_array_muxed2;
			end
			7'd84: begin
				storav84 <= sync_array_muxed2;
			end
			7'd85: begin
				storav85 <= sync_array_muxed2;
			end
			7'd86: begin
				storav86 <= sync_array_muxed2;
			end
			7'd87: begin
				storav87 <= sync_array_muxed2;
			end
			7'd88: begin
				storav88 <= sync_array_muxed2;
			end
			7'd89: begin
				storav89 <= sync_array_muxed2;
			end
			7'd90: begin
				storav90 <= sync_array_muxed2;
			end
			7'd91: begin
				storav91 <= sync_array_muxed2;
			end
			7'd92: begin
				storav92 <= sync_array_muxed2;
			end
			7'd93: begin
				storav93 <= sync_array_muxed2;
			end
			7'd94: begin
				storav94 <= sync_array_muxed2;
			end
			7'd95: begin
				storav95 <= sync_array_muxed2;
			end
			7'd96: begin
				storav96 <= sync_array_muxed2;
			end
			7'd97: begin
				storav97 <= sync_array_muxed2;
			end
			7'd98: begin
				storav98 <= sync_array_muxed2;
			end
			7'd99: begin
				storav99 <= sync_array_muxed2;
			end
			7'd100: begin
				storav100 <= sync_array_muxed2;
			end
			7'd101: begin
				storav101 <= sync_array_muxed2;
			end
			7'd102: begin
				storav102 <= sync_array_muxed2;
			end
			7'd103: begin
				storav103 <= sync_array_muxed2;
			end
			7'd104: begin
				storav104 <= sync_array_muxed2;
			end
			7'd105: begin
				storav105 <= sync_array_muxed2;
			end
			7'd106: begin
				storav106 <= sync_array_muxed2;
			end
			7'd107: begin
				storav107 <= sync_array_muxed2;
			end
			7'd108: begin
				storav108 <= sync_array_muxed2;
			end
			7'd109: begin
				storav109 <= sync_array_muxed2;
			end
			7'd110: begin
				storav110 <= sync_array_muxed2;
			end
			7'd111: begin
				storav111 <= sync_array_muxed2;
			end
			7'd112: begin
				storav112 <= sync_array_muxed2;
			end
			7'd113: begin
				storav113 <= sync_array_muxed2;
			end
			7'd114: begin
				storav114 <= sync_array_muxed2;
			end
			7'd115: begin
				storav115 <= sync_array_muxed2;
			end
			7'd116: begin
				storav116 <= sync_array_muxed2;
			end
			7'd117: begin
				storav117 <= sync_array_muxed2;
			end
			7'd118: begin
				storav118 <= sync_array_muxed2;
			end
			7'd119: begin
				storav119 <= sync_array_muxed2;
			end
			7'd120: begin
				storav120 <= sync_array_muxed2;
			end
			7'd121: begin
				storav121 <= sync_array_muxed2;
			end
			7'd122: begin
				storav122 <= sync_array_muxed2;
			end
			7'd123: begin
				storav123 <= sync_array_muxed2;
			end
			7'd124: begin
				storav124 <= sync_array_muxed2;
			end
			7'd125: begin
				storav125 <= sync_array_muxed2;
			end
			7'd126: begin
				storav126 <= sync_array_muxed2;
			end
			default: begin
				storav127 <= sync_array_muxed2;
			end
		endcase
	end
	if (f_next_value_ce1) begin
		sync_array_muxed3 = f_next_value1;
		case (ADR_i)
			1'd0: begin
				storak0 <= sync_array_muxed3;
			end
			1'd1: begin
				storak1 <= sync_array_muxed3;
			end
			2'd2: begin
				storak2 <= sync_array_muxed3;
			end
			2'd3: begin
				storak3 <= sync_array_muxed3;
			end
			3'd4: begin
				storak4 <= sync_array_muxed3;
			end
			3'd5: begin
				storak5 <= sync_array_muxed3;
			end
			3'd6: begin
				storak6 <= sync_array_muxed3;
			end
			3'd7: begin
				storak7 <= sync_array_muxed3;
			end
			4'd8: begin
				storak8 <= sync_array_muxed3;
			end
			4'd9: begin
				storak9 <= sync_array_muxed3;
			end
			4'd10: begin
				storak10 <= sync_array_muxed3;
			end
			4'd11: begin
				storak11 <= sync_array_muxed3;
			end
			4'd12: begin
				storak12 <= sync_array_muxed3;
			end
			4'd13: begin
				storak13 <= sync_array_muxed3;
			end
			4'd14: begin
				storak14 <= sync_array_muxed3;
			end
			4'd15: begin
				storak15 <= sync_array_muxed3;
			end
			5'd16: begin
				storak16 <= sync_array_muxed3;
			end
			5'd17: begin
				storak17 <= sync_array_muxed3;
			end
			5'd18: begin
				storak18 <= sync_array_muxed3;
			end
			5'd19: begin
				storak19 <= sync_array_muxed3;
			end
			5'd20: begin
				storak20 <= sync_array_muxed3;
			end
			5'd21: begin
				storak21 <= sync_array_muxed3;
			end
			5'd22: begin
				storak22 <= sync_array_muxed3;
			end
			5'd23: begin
				storak23 <= sync_array_muxed3;
			end
			5'd24: begin
				storak24 <= sync_array_muxed3;
			end
			5'd25: begin
				storak25 <= sync_array_muxed3;
			end
			5'd26: begin
				storak26 <= sync_array_muxed3;
			end
			5'd27: begin
				storak27 <= sync_array_muxed3;
			end
			5'd28: begin
				storak28 <= sync_array_muxed3;
			end
			5'd29: begin
				storak29 <= sync_array_muxed3;
			end
			5'd30: begin
				storak30 <= sync_array_muxed3;
			end
			5'd31: begin
				storak31 <= sync_array_muxed3;
			end
			6'd32: begin
				storak32 <= sync_array_muxed3;
			end
			6'd33: begin
				storak33 <= sync_array_muxed3;
			end
			6'd34: begin
				storak34 <= sync_array_muxed3;
			end
			6'd35: begin
				storak35 <= sync_array_muxed3;
			end
			6'd36: begin
				storak36 <= sync_array_muxed3;
			end
			6'd37: begin
				storak37 <= sync_array_muxed3;
			end
			6'd38: begin
				storak38 <= sync_array_muxed3;
			end
			6'd39: begin
				storak39 <= sync_array_muxed3;
			end
			6'd40: begin
				storak40 <= sync_array_muxed3;
			end
			6'd41: begin
				storak41 <= sync_array_muxed3;
			end
			6'd42: begin
				storak42 <= sync_array_muxed3;
			end
			6'd43: begin
				storak43 <= sync_array_muxed3;
			end
			6'd44: begin
				storak44 <= sync_array_muxed3;
			end
			6'd45: begin
				storak45 <= sync_array_muxed3;
			end
			6'd46: begin
				storak46 <= sync_array_muxed3;
			end
			6'd47: begin
				storak47 <= sync_array_muxed3;
			end
			6'd48: begin
				storak48 <= sync_array_muxed3;
			end
			6'd49: begin
				storak49 <= sync_array_muxed3;
			end
			6'd50: begin
				storak50 <= sync_array_muxed3;
			end
			6'd51: begin
				storak51 <= sync_array_muxed3;
			end
			6'd52: begin
				storak52 <= sync_array_muxed3;
			end
			6'd53: begin
				storak53 <= sync_array_muxed3;
			end
			6'd54: begin
				storak54 <= sync_array_muxed3;
			end
			6'd55: begin
				storak55 <= sync_array_muxed3;
			end
			6'd56: begin
				storak56 <= sync_array_muxed3;
			end
			6'd57: begin
				storak57 <= sync_array_muxed3;
			end
			6'd58: begin
				storak58 <= sync_array_muxed3;
			end
			6'd59: begin
				storak59 <= sync_array_muxed3;
			end
			6'd60: begin
				storak60 <= sync_array_muxed3;
			end
			6'd61: begin
				storak61 <= sync_array_muxed3;
			end
			6'd62: begin
				storak62 <= sync_array_muxed3;
			end
			6'd63: begin
				storak63 <= sync_array_muxed3;
			end
			7'd64: begin
				storak64 <= sync_array_muxed3;
			end
			7'd65: begin
				storak65 <= sync_array_muxed3;
			end
			7'd66: begin
				storak66 <= sync_array_muxed3;
			end
			7'd67: begin
				storak67 <= sync_array_muxed3;
			end
			7'd68: begin
				storak68 <= sync_array_muxed3;
			end
			7'd69: begin
				storak69 <= sync_array_muxed3;
			end
			7'd70: begin
				storak70 <= sync_array_muxed3;
			end
			7'd71: begin
				storak71 <= sync_array_muxed3;
			end
			7'd72: begin
				storak72 <= sync_array_muxed3;
			end
			7'd73: begin
				storak73 <= sync_array_muxed3;
			end
			7'd74: begin
				storak74 <= sync_array_muxed3;
			end
			7'd75: begin
				storak75 <= sync_array_muxed3;
			end
			7'd76: begin
				storak76 <= sync_array_muxed3;
			end
			7'd77: begin
				storak77 <= sync_array_muxed3;
			end
			7'd78: begin
				storak78 <= sync_array_muxed3;
			end
			7'd79: begin
				storak79 <= sync_array_muxed3;
			end
			7'd80: begin
				storak80 <= sync_array_muxed3;
			end
			7'd81: begin
				storak81 <= sync_array_muxed3;
			end
			7'd82: begin
				storak82 <= sync_array_muxed3;
			end
			7'd83: begin
				storak83 <= sync_array_muxed3;
			end
			7'd84: begin
				storak84 <= sync_array_muxed3;
			end
			7'd85: begin
				storak85 <= sync_array_muxed3;
			end
			7'd86: begin
				storak86 <= sync_array_muxed3;
			end
			7'd87: begin
				storak87 <= sync_array_muxed3;
			end
			7'd88: begin
				storak88 <= sync_array_muxed3;
			end
			7'd89: begin
				storak89 <= sync_array_muxed3;
			end
			7'd90: begin
				storak90 <= sync_array_muxed3;
			end
			7'd91: begin
				storak91 <= sync_array_muxed3;
			end
			7'd92: begin
				storak92 <= sync_array_muxed3;
			end
			7'd93: begin
				storak93 <= sync_array_muxed3;
			end
			7'd94: begin
				storak94 <= sync_array_muxed3;
			end
			7'd95: begin
				storak95 <= sync_array_muxed3;
			end
			7'd96: begin
				storak96 <= sync_array_muxed3;
			end
			7'd97: begin
				storak97 <= sync_array_muxed3;
			end
			7'd98: begin
				storak98 <= sync_array_muxed3;
			end
			7'd99: begin
				storak99 <= sync_array_muxed3;
			end
			7'd100: begin
				storak100 <= sync_array_muxed3;
			end
			7'd101: begin
				storak101 <= sync_array_muxed3;
			end
			7'd102: begin
				storak102 <= sync_array_muxed3;
			end
			7'd103: begin
				storak103 <= sync_array_muxed3;
			end
			7'd104: begin
				storak104 <= sync_array_muxed3;
			end
			7'd105: begin
				storak105 <= sync_array_muxed3;
			end
			7'd106: begin
				storak106 <= sync_array_muxed3;
			end
			7'd107: begin
				storak107 <= sync_array_muxed3;
			end
			7'd108: begin
				storak108 <= sync_array_muxed3;
			end
			7'd109: begin
				storak109 <= sync_array_muxed3;
			end
			7'd110: begin
				storak110 <= sync_array_muxed3;
			end
			7'd111: begin
				storak111 <= sync_array_muxed3;
			end
			7'd112: begin
				storak112 <= sync_array_muxed3;
			end
			7'd113: begin
				storak113 <= sync_array_muxed3;
			end
			7'd114: begin
				storak114 <= sync_array_muxed3;
			end
			7'd115: begin
				storak115 <= sync_array_muxed3;
			end
			7'd116: begin
				storak116 <= sync_array_muxed3;
			end
			7'd117: begin
				storak117 <= sync_array_muxed3;
			end
			7'd118: begin
				storak118 <= sync_array_muxed3;
			end
			7'd119: begin
				storak119 <= sync_array_muxed3;
			end
			7'd120: begin
				storak120 <= sync_array_muxed3;
			end
			7'd121: begin
				storak121 <= sync_array_muxed3;
			end
			7'd122: begin
				storak122 <= sync_array_muxed3;
			end
			7'd123: begin
				storak123 <= sync_array_muxed3;
			end
			7'd124: begin
				storak124 <= sync_array_muxed3;
			end
			7'd125: begin
				storak125 <= sync_array_muxed3;
			end
			7'd126: begin
				storak126 <= sync_array_muxed3;
			end
			default: begin
				storak127 <= sync_array_muxed3;
			end
		endcase
	end
	if (sys_rst) begin
		STALL_o <= 1'd0;
		ACK_o <= 1'd0;
		DAT_o <= 64'd0;
		storak0 <= 64'd0;
		storak1 <= 64'd0;
		storak2 <= 64'd0;
		storak3 <= 64'd0;
		storak4 <= 64'd0;
		storak5 <= 64'd0;
		storak6 <= 64'd0;
		storak7 <= 64'd0;
		storak8 <= 64'd0;
		storak9 <= 64'd0;
		storak10 <= 64'd0;
		storak11 <= 64'd0;
		storak12 <= 64'd0;
		storak13 <= 64'd0;
		storak14 <= 64'd0;
		storak15 <= 64'd0;
		storak16 <= 64'd0;
		storak17 <= 64'd0;
		storak18 <= 64'd0;
		storak19 <= 64'd0;
		storak20 <= 64'd0;
		storak21 <= 64'd0;
		storak22 <= 64'd0;
		storak23 <= 64'd0;
		storak24 <= 64'd0;
		storak25 <= 64'd0;
		storak26 <= 64'd0;
		storak27 <= 64'd0;
		storak28 <= 64'd0;
		storak29 <= 64'd0;
		storak30 <= 64'd0;
		storak31 <= 64'd0;
		storak32 <= 64'd0;
		storak33 <= 64'd0;
		storak34 <= 64'd0;
		storak35 <= 64'd0;
		storak36 <= 64'd0;
		storak37 <= 64'd0;
		storak38 <= 64'd0;
		storak39 <= 64'd0;
		storak40 <= 64'd0;
		storak41 <= 64'd0;
		storak42 <= 64'd0;
		storak43 <= 64'd0;
		storak44 <= 64'd0;
		storak45 <= 64'd0;
		storak46 <= 64'd0;
		storak47 <= 64'd0;
		storak48 <= 64'd0;
		storak49 <= 64'd0;
		storak50 <= 64'd0;
		storak51 <= 64'd0;
		storak52 <= 64'd0;
		storak53 <= 64'd0;
		storak54 <= 64'd0;
		storak55 <= 64'd0;
		storak56 <= 64'd0;
		storak57 <= 64'd0;
		storak58 <= 64'd0;
		storak59 <= 64'd0;
		storak60 <= 64'd0;
		storak61 <= 64'd0;
		storak62 <= 64'd0;
		storak63 <= 64'd0;
		storak64 <= 64'd0;
		storak65 <= 64'd0;
		storak66 <= 64'd0;
		storak67 <= 64'd0;
		storak68 <= 64'd0;
		storak69 <= 64'd0;
		storak70 <= 64'd0;
		storak71 <= 64'd0;
		storak72 <= 64'd0;
		storak73 <= 64'd0;
		storak74 <= 64'd0;
		storak75 <= 64'd0;
		storak76 <= 64'd0;
		storak77 <= 64'd0;
		storak78 <= 64'd0;
		storak79 <= 64'd0;
		storak80 <= 64'd0;
		storak81 <= 64'd0;
		storak82 <= 64'd0;
		storak83 <= 64'd0;
		storak84 <= 64'd0;
		storak85 <= 64'd0;
		storak86 <= 64'd0;
		storak87 <= 64'd0;
		storak88 <= 64'd0;
		storak89 <= 64'd0;
		storak90 <= 64'd0;
		storak91 <= 64'd0;
		storak92 <= 64'd0;
		storak93 <= 64'd0;
		storak94 <= 64'd0;
		storak95 <= 64'd0;
		storak96 <= 64'd0;
		storak97 <= 64'd0;
		storak98 <= 64'd0;
		storak99 <= 64'd0;
		storak100 <= 64'd0;
		storak101 <= 64'd0;
		storak102 <= 64'd0;
		storak103 <= 64'd0;
		storak104 <= 64'd0;
		storak105 <= 64'd0;
		storak106 <= 64'd0;
		storak107 <= 64'd0;
		storak108 <= 64'd0;
		storak109 <= 64'd0;
		storak110 <= 64'd0;
		storak111 <= 64'd0;
		storak112 <= 64'd0;
		storak113 <= 64'd0;
		storak114 <= 64'd0;
		storak115 <= 64'd0;
		storak116 <= 64'd0;
		storak117 <= 64'd0;
		storak118 <= 64'd0;
		storak119 <= 64'd0;
		storak120 <= 64'd0;
		storak121 <= 64'd0;
		storak122 <= 64'd0;
		storak123 <= 64'd0;
		storak124 <= 64'd0;
		storak125 <= 64'd0;
		storak126 <= 64'd0;
		storak127 <= 64'd0;
		storav0 <= 64'd0;
		storav1 <= 64'd0;
		storav2 <= 64'd0;
		storav3 <= 64'd0;
		storav4 <= 64'd0;
		storav5 <= 64'd0;
		storav6 <= 64'd0;
		storav7 <= 64'd0;
		storav8 <= 64'd0;
		storav9 <= 64'd0;
		storav10 <= 64'd0;
		storav11 <= 64'd0;
		storav12 <= 64'd0;
		storav13 <= 64'd0;
		storav14 <= 64'd0;
		storav15 <= 64'd0;
		storav16 <= 64'd0;
		storav17 <= 64'd0;
		storav18 <= 64'd0;
		storav19 <= 64'd0;
		storav20 <= 64'd0;
		storav21 <= 64'd0;
		storav22 <= 64'd0;
		storav23 <= 64'd0;
		storav24 <= 64'd0;
		storav25 <= 64'd0;
		storav26 <= 64'd0;
		storav27 <= 64'd0;
		storav28 <= 64'd0;
		storav29 <= 64'd0;
		storav30 <= 64'd0;
		storav31 <= 64'd0;
		storav32 <= 64'd0;
		storav33 <= 64'd0;
		storav34 <= 64'd0;
		storav35 <= 64'd0;
		storav36 <= 64'd0;
		storav37 <= 64'd0;
		storav38 <= 64'd0;
		storav39 <= 64'd0;
		storav40 <= 64'd0;
		storav41 <= 64'd0;
		storav42 <= 64'd0;
		storav43 <= 64'd0;
		storav44 <= 64'd0;
		storav45 <= 64'd0;
		storav46 <= 64'd0;
		storav47 <= 64'd0;
		storav48 <= 64'd0;
		storav49 <= 64'd0;
		storav50 <= 64'd0;
		storav51 <= 64'd0;
		storav52 <= 64'd0;
		storav53 <= 64'd0;
		storav54 <= 64'd0;
		storav55 <= 64'd0;
		storav56 <= 64'd0;
		storav57 <= 64'd0;
		storav58 <= 64'd0;
		storav59 <= 64'd0;
		storav60 <= 64'd0;
		storav61 <= 64'd0;
		storav62 <= 64'd0;
		storav63 <= 64'd0;
		storav64 <= 64'd0;
		storav65 <= 64'd0;
		storav66 <= 64'd0;
		storav67 <= 64'd0;
		storav68 <= 64'd0;
		storav69 <= 64'd0;
		storav70 <= 64'd0;
		storav71 <= 64'd0;
		storav72 <= 64'd0;
		storav73 <= 64'd0;
		storav74 <= 64'd0;
		storav75 <= 64'd0;
		storav76 <= 64'd0;
		storav77 <= 64'd0;
		storav78 <= 64'd0;
		storav79 <= 64'd0;
		storav80 <= 64'd0;
		storav81 <= 64'd0;
		storav82 <= 64'd0;
		storav83 <= 64'd0;
		storav84 <= 64'd0;
		storav85 <= 64'd0;
		storav86 <= 64'd0;
		storav87 <= 64'd0;
		storav88 <= 64'd0;
		storav89 <= 64'd0;
		storav90 <= 64'd0;
		storav91 <= 64'd0;
		storav92 <= 64'd0;
		storav93 <= 64'd0;
		storav94 <= 64'd0;
		storav95 <= 64'd0;
		storav96 <= 64'd0;
		storav97 <= 64'd0;
		storav98 <= 64'd0;
		storav99 <= 64'd0;
		storav100 <= 64'd0;
		storav101 <= 64'd0;
		storav102 <= 64'd0;
		storav103 <= 64'd0;
		storav104 <= 64'd0;
		storav105 <= 64'd0;
		storav106 <= 64'd0;
		storav107 <= 64'd0;
		storav108 <= 64'd0;
		storav109 <= 64'd0;
		storav110 <= 64'd0;
		storav111 <= 64'd0;
		storav112 <= 64'd0;
		storav113 <= 64'd0;
		storav114 <= 64'd0;
		storav115 <= 64'd0;
		storav116 <= 64'd0;
		storav117 <= 64'd0;
		storav118 <= 64'd0;
		storav119 <= 64'd0;
		storav120 <= 64'd0;
		storav121 <= 64'd0;
		storav122 <= 64'd0;
		storav123 <= 64'd0;
		storav124 <= 64'd0;
		storav125 <= 64'd0;
		storav126 <= 64'd0;
		storav127 <= 64'd0;
		empty_location <= 64'd0;
		state <= 2'd3;
	end
end

endmodule


