/* Machine-generated using Migen */
module keyvalue_3(
	input sys_rst,
	input [3:0] SEL_i,
	input ADR_IS_KEY_i,
	input DAT_IS_KEY_i,
	input [15:0] ADR_i,
	input [15:0] DAT_i,
	input WE_i,
	input STB_i,
	input CYC_i,
	output reg DUP_o,
	output reg STALL_o,
	output reg ACK_o,
	output reg [15:0] DAT_o,
	output [15:0] LA_o,
	input sys_clk,
	input sys_rst_1
);

reg [15:0] __main___storak0 = 16'd0;
reg [15:0] __main___storak1 = 16'd0;
reg [15:0] __main___storak2 = 16'd0;
reg [15:0] __main___storak3 = 16'd0;
reg [15:0] __main___storak4 = 16'd0;
reg [15:0] __main___storak5 = 16'd0;
reg [15:0] __main___storak6 = 16'd0;
reg [15:0] __main___storak7 = 16'd0;
reg [15:0] __main___storak8 = 16'd0;
reg [15:0] __main___storak9 = 16'd0;
reg [15:0] __main___storak10 = 16'd0;
reg [15:0] __main___storak11 = 16'd0;
reg [15:0] __main___storak12 = 16'd0;
reg [15:0] __main___storak13 = 16'd0;
reg [15:0] __main___storak14 = 16'd0;
reg [15:0] __main___storak15 = 16'd0;
reg [15:0] __main___storak16 = 16'd0;
reg [15:0] __main___storak17 = 16'd0;
reg [15:0] __main___storak18 = 16'd0;
reg [15:0] __main___storak19 = 16'd0;
reg [15:0] __main___storak20 = 16'd0;
reg [15:0] __main___storak21 = 16'd0;
reg [15:0] __main___storak22 = 16'd0;
reg [15:0] __main___storak23 = 16'd0;
reg [15:0] __main___storak24 = 16'd0;
reg [15:0] __main___storak25 = 16'd0;
reg [15:0] __main___storak26 = 16'd0;
reg [15:0] __main___storak27 = 16'd0;
reg [15:0] __main___storak28 = 16'd0;
reg [15:0] __main___storak29 = 16'd0;
reg [15:0] __main___storak30 = 16'd0;
reg [15:0] __main___storak31 = 16'd0;
reg [15:0] __main___storav0 = 16'd0;
reg [15:0] __main___storav1 = 16'd0;
reg [15:0] __main___storav2 = 16'd0;
reg [15:0] __main___storav3 = 16'd0;
reg [15:0] __main___storav4 = 16'd0;
reg [15:0] __main___storav5 = 16'd0;
reg [15:0] __main___storav6 = 16'd0;
reg [15:0] __main___storav7 = 16'd0;
reg [15:0] __main___storav8 = 16'd0;
reg [15:0] __main___storav9 = 16'd0;
reg [15:0] __main___storav10 = 16'd0;
reg [15:0] __main___storav11 = 16'd0;
reg [15:0] __main___storav12 = 16'd0;
reg [15:0] __main___storav13 = 16'd0;
reg [15:0] __main___storav14 = 16'd0;
reg [15:0] __main___storav15 = 16'd0;
reg [15:0] __main___storav16 = 16'd0;
reg [15:0] __main___storav17 = 16'd0;
reg [15:0] __main___storav18 = 16'd0;
reg [15:0] __main___storav19 = 16'd0;
reg [15:0] __main___storav20 = 16'd0;
reg [15:0] __main___storav21 = 16'd0;
reg [15:0] __main___storav22 = 16'd0;
reg [15:0] __main___storav23 = 16'd0;
reg [15:0] __main___storav24 = 16'd0;
reg [15:0] __main___storav25 = 16'd0;
reg [15:0] __main___storav26 = 16'd0;
reg [15:0] __main___storav27 = 16'd0;
reg [15:0] __main___storav28 = 16'd0;
reg [15:0] __main___storav29 = 16'd0;
reg [15:0] __main___storav30 = 16'd0;
reg [15:0] __main___storav31 = 16'd0;
reg [15:0] __main___empty_location = 16'd1;
reg [1:0] convert_state = 2'd3;
reg [1:0] convert_next_state;
reg __main___STALL_o_next_value0;
reg __main___STALL_o_next_value_ce0;
reg [15:0] __main___empty_location_t_next_value;
reg __main___empty_location_t_next_value_ce;
reg __main___ACK_o_f_next_value;
reg __main___ACK_o_f_next_value_ce;
reg [15:0] __main___DAT_o_next_value1;
reg __main___DAT_o_next_value_ce1;
reg __main___DUP_o_next_value2;
reg __main___DUP_o_next_value_ce2;
reg [15:0] convert_next_value0;
reg convert_next_value_ce0;
reg [15:0] convert_next_value1;
reg convert_next_value_ce1;
reg [15:0] convert_t_next_value;
reg convert_t_next_value_ce;
reg [15:0] convert_f_next_value;
reg convert_f_next_value_ce;
reg [15:0] convert_comb_array_muxed;
reg [15:0] convert_sync_array_muxed0 = 16'd0;
reg [15:0] convert_sync_array_muxed1 = 16'd0;
reg [15:0] convert_sync_array_muxed2 = 16'd0;
reg [15:0] convert_sync_array_muxed3 = 16'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign LA_o = DAT_o;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	convert_next_state <= 2'd0;
	__main___STALL_o_next_value0 <= 1'd0;
	__main___STALL_o_next_value_ce0 <= 1'd0;
	__main___empty_location_t_next_value <= 16'd0;
	__main___empty_location_t_next_value_ce <= 1'd0;
	__main___ACK_o_f_next_value <= 1'd0;
	__main___ACK_o_f_next_value_ce <= 1'd0;
	__main___DAT_o_next_value1 <= 16'd0;
	__main___DAT_o_next_value_ce1 <= 1'd0;
	__main___DUP_o_next_value2 <= 1'd0;
	__main___DUP_o_next_value_ce2 <= 1'd0;
	convert_next_value0 <= 16'd0;
	convert_next_value_ce0 <= 1'd0;
	convert_next_value1 <= 16'd0;
	convert_next_value_ce1 <= 1'd0;
	convert_t_next_value <= 16'd0;
	convert_t_next_value_ce <= 1'd0;
	convert_f_next_value <= 16'd0;
	convert_f_next_value_ce <= 1'd0;
	convert_next_state <= convert_state;
	case (convert_state)
		1'd0: begin
			__main___STALL_o_next_value0 <= 1'd0;
			__main___STALL_o_next_value_ce0 <= 1'd1;
			if ((((STB_i == 1'd1) & (WE_i == 1'd0)) & (ACK_o == 1'd0))) begin
				convert_next_state <= 1'd1;
			end else begin
				if ((((STB_i == 1'd1) & (WE_i == 1'd1)) & (ACK_o == 1'd0))) begin
					convert_next_state <= 2'd2;
					if (ADR_IS_KEY_i) begin
						__main___empty_location_t_next_value <= (__main___empty_location + 1'd1);
						__main___empty_location_t_next_value_ce <= 1'd1;
					end
				end else begin
					__main___ACK_o_f_next_value <= 1'd0;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
		end
		1'd1: begin
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak1 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav1;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav1 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak1;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak2 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav2;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav2 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak2;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak3 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav3;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav3 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak3;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak4 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav4;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav4 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak4;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak5 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav5;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav5 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak5;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak6 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav6;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav6 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak6;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak7 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav7;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav7 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak7;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak8 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav8;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav8 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak8;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak9 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav9;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav9 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak9;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak10 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav10;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav10 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak10;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak11 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav11;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav11 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak11;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak12 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav12;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav12 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak12;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak13 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav13;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav13 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak13;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak14 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav14;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav14 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak14;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak15 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav15;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav15 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak15;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak16 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav16;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav16 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak16;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak17 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav17;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav17 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak17;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak18 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav18;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav18 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak18;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak19 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav19;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav19 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak19;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak20 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav20;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav20 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak20;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak21 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav21;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav21 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak21;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak22 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav22;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav22 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak22;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak23 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav23;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav23 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak23;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak24 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav24;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav24 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak24;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak25 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav25;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav25 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak25;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak26 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav26;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav26 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak26;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak27 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav27;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav27 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak27;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak28 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav28;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav28 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak28;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak29 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav29;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav29 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak29;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak30 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav30;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav30 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak30;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak31 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav31;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((DAT_i > 1'd0)) begin
				if ((__main___storav31 == DAT_i)) begin
					__main___DAT_o_next_value1 <= __main___storak31;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd0)) begin
				if ((ADR_i == 1'd0)) begin
					if ((DAT_i == 1'd0)) begin
						__main___ACK_o_f_next_value <= 1'd1;
						__main___ACK_o_f_next_value_ce <= 1'd1;
						__main___DUP_o_next_value2 <= 1'd1;
						__main___DUP_o_next_value_ce2 <= 1'd1;
						__main___DAT_o_next_value1 <= 1'sd1;
						__main___DAT_o_next_value_ce1 <= 1'd1;
					end
				end else begin
					__main___DAT_o_next_value1 <= convert_comb_array_muxed;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((sys_rst == 1'd1)) begin
				convert_next_state <= 2'd3;
			end
		end
		2'd2: begin
			if (ADR_IS_KEY_i) begin
				convert_next_value0 <= DAT_i;
				convert_next_value_ce0 <= 1'd1;
				convert_next_value1 <= ADR_i;
				convert_next_value_ce1 <= 1'd1;
				__main___DAT_o_next_value1 <= __main___empty_location;
				__main___DAT_o_next_value_ce1 <= 1'd1;
			end else begin
				if (DAT_IS_KEY_i) begin
					convert_t_next_value <= DAT_i;
					convert_t_next_value_ce <= 1'd1;
					__main___DAT_o_next_value1 <= ADR_i;
					__main___DAT_o_next_value_ce1 <= 1'd1;
				end else begin
					convert_f_next_value <= DAT_i;
					convert_f_next_value_ce <= 1'd1;
					__main___DAT_o_next_value1 <= ADR_i;
					__main___DAT_o_next_value_ce1 <= 1'd1;
				end
			end
			__main___ACK_o_f_next_value <= 1'd1;
			__main___ACK_o_f_next_value_ce <= 1'd1;
			convert_next_state <= 1'd0;
			if ((sys_rst == 1'd1)) begin
				convert_next_state <= 2'd3;
			end else begin
				convert_next_state <= 1'd0;
			end
		end
		default: begin
			convert_next_state <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	convert_comb_array_muxed <= 16'd0;
	case (ADR_i)
		1'd0: begin
			convert_comb_array_muxed <= __main___storav0;
		end
		1'd1: begin
			convert_comb_array_muxed <= __main___storav1;
		end
		2'd2: begin
			convert_comb_array_muxed <= __main___storav2;
		end
		2'd3: begin
			convert_comb_array_muxed <= __main___storav3;
		end
		3'd4: begin
			convert_comb_array_muxed <= __main___storav4;
		end
		3'd5: begin
			convert_comb_array_muxed <= __main___storav5;
		end
		3'd6: begin
			convert_comb_array_muxed <= __main___storav6;
		end
		3'd7: begin
			convert_comb_array_muxed <= __main___storav7;
		end
		4'd8: begin
			convert_comb_array_muxed <= __main___storav8;
		end
		4'd9: begin
			convert_comb_array_muxed <= __main___storav9;
		end
		4'd10: begin
			convert_comb_array_muxed <= __main___storav10;
		end
		4'd11: begin
			convert_comb_array_muxed <= __main___storav11;
		end
		4'd12: begin
			convert_comb_array_muxed <= __main___storav12;
		end
		4'd13: begin
			convert_comb_array_muxed <= __main___storav13;
		end
		4'd14: begin
			convert_comb_array_muxed <= __main___storav14;
		end
		4'd15: begin
			convert_comb_array_muxed <= __main___storav15;
		end
		5'd16: begin
			convert_comb_array_muxed <= __main___storav16;
		end
		5'd17: begin
			convert_comb_array_muxed <= __main___storav17;
		end
		5'd18: begin
			convert_comb_array_muxed <= __main___storav18;
		end
		5'd19: begin
			convert_comb_array_muxed <= __main___storav19;
		end
		5'd20: begin
			convert_comb_array_muxed <= __main___storav20;
		end
		5'd21: begin
			convert_comb_array_muxed <= __main___storav21;
		end
		5'd22: begin
			convert_comb_array_muxed <= __main___storav22;
		end
		5'd23: begin
			convert_comb_array_muxed <= __main___storav23;
		end
		5'd24: begin
			convert_comb_array_muxed <= __main___storav24;
		end
		5'd25: begin
			convert_comb_array_muxed <= __main___storav25;
		end
		5'd26: begin
			convert_comb_array_muxed <= __main___storav26;
		end
		5'd27: begin
			convert_comb_array_muxed <= __main___storav27;
		end
		5'd28: begin
			convert_comb_array_muxed <= __main___storav28;
		end
		5'd29: begin
			convert_comb_array_muxed <= __main___storav29;
		end
		5'd30: begin
			convert_comb_array_muxed <= __main___storav30;
		end
		default: begin
			convert_comb_array_muxed <= __main___storav31;
		end
	endcase
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

always @(posedge sys_clk) begin
	convert_state <= convert_next_state;
	if (__main___STALL_o_next_value_ce0) begin
		STALL_o <= __main___STALL_o_next_value0;
	end
	if (__main___empty_location_t_next_value_ce) begin
		__main___empty_location <= __main___empty_location_t_next_value;
	end
	if (__main___ACK_o_f_next_value_ce) begin
		ACK_o <= __main___ACK_o_f_next_value;
	end
	if (__main___DAT_o_next_value_ce1) begin
		DAT_o <= __main___DAT_o_next_value1;
	end
	if (__main___DUP_o_next_value_ce2) begin
		DUP_o <= __main___DUP_o_next_value2;
	end
	if (convert_next_value_ce0) begin
		convert_sync_array_muxed0 = convert_next_value0;
		case (__main___empty_location)
			1'd0: begin
				__main___storav0 <= convert_sync_array_muxed0;
			end
			1'd1: begin
				__main___storav1 <= convert_sync_array_muxed0;
			end
			2'd2: begin
				__main___storav2 <= convert_sync_array_muxed0;
			end
			2'd3: begin
				__main___storav3 <= convert_sync_array_muxed0;
			end
			3'd4: begin
				__main___storav4 <= convert_sync_array_muxed0;
			end
			3'd5: begin
				__main___storav5 <= convert_sync_array_muxed0;
			end
			3'd6: begin
				__main___storav6 <= convert_sync_array_muxed0;
			end
			3'd7: begin
				__main___storav7 <= convert_sync_array_muxed0;
			end
			4'd8: begin
				__main___storav8 <= convert_sync_array_muxed0;
			end
			4'd9: begin
				__main___storav9 <= convert_sync_array_muxed0;
			end
			4'd10: begin
				__main___storav10 <= convert_sync_array_muxed0;
			end
			4'd11: begin
				__main___storav11 <= convert_sync_array_muxed0;
			end
			4'd12: begin
				__main___storav12 <= convert_sync_array_muxed0;
			end
			4'd13: begin
				__main___storav13 <= convert_sync_array_muxed0;
			end
			4'd14: begin
				__main___storav14 <= convert_sync_array_muxed0;
			end
			4'd15: begin
				__main___storav15 <= convert_sync_array_muxed0;
			end
			5'd16: begin
				__main___storav16 <= convert_sync_array_muxed0;
			end
			5'd17: begin
				__main___storav17 <= convert_sync_array_muxed0;
			end
			5'd18: begin
				__main___storav18 <= convert_sync_array_muxed0;
			end
			5'd19: begin
				__main___storav19 <= convert_sync_array_muxed0;
			end
			5'd20: begin
				__main___storav20 <= convert_sync_array_muxed0;
			end
			5'd21: begin
				__main___storav21 <= convert_sync_array_muxed0;
			end
			5'd22: begin
				__main___storav22 <= convert_sync_array_muxed0;
			end
			5'd23: begin
				__main___storav23 <= convert_sync_array_muxed0;
			end
			5'd24: begin
				__main___storav24 <= convert_sync_array_muxed0;
			end
			5'd25: begin
				__main___storav25 <= convert_sync_array_muxed0;
			end
			5'd26: begin
				__main___storav26 <= convert_sync_array_muxed0;
			end
			5'd27: begin
				__main___storav27 <= convert_sync_array_muxed0;
			end
			5'd28: begin
				__main___storav28 <= convert_sync_array_muxed0;
			end
			5'd29: begin
				__main___storav29 <= convert_sync_array_muxed0;
			end
			5'd30: begin
				__main___storav30 <= convert_sync_array_muxed0;
			end
			default: begin
				__main___storav31 <= convert_sync_array_muxed0;
			end
		endcase
	end
	if (convert_next_value_ce1) begin
		convert_sync_array_muxed1 = convert_next_value1;
		case (__main___empty_location)
			1'd0: begin
				__main___storak0 <= convert_sync_array_muxed1;
			end
			1'd1: begin
				__main___storak1 <= convert_sync_array_muxed1;
			end
			2'd2: begin
				__main___storak2 <= convert_sync_array_muxed1;
			end
			2'd3: begin
				__main___storak3 <= convert_sync_array_muxed1;
			end
			3'd4: begin
				__main___storak4 <= convert_sync_array_muxed1;
			end
			3'd5: begin
				__main___storak5 <= convert_sync_array_muxed1;
			end
			3'd6: begin
				__main___storak6 <= convert_sync_array_muxed1;
			end
			3'd7: begin
				__main___storak7 <= convert_sync_array_muxed1;
			end
			4'd8: begin
				__main___storak8 <= convert_sync_array_muxed1;
			end
			4'd9: begin
				__main___storak9 <= convert_sync_array_muxed1;
			end
			4'd10: begin
				__main___storak10 <= convert_sync_array_muxed1;
			end
			4'd11: begin
				__main___storak11 <= convert_sync_array_muxed1;
			end
			4'd12: begin
				__main___storak12 <= convert_sync_array_muxed1;
			end
			4'd13: begin
				__main___storak13 <= convert_sync_array_muxed1;
			end
			4'd14: begin
				__main___storak14 <= convert_sync_array_muxed1;
			end
			4'd15: begin
				__main___storak15 <= convert_sync_array_muxed1;
			end
			5'd16: begin
				__main___storak16 <= convert_sync_array_muxed1;
			end
			5'd17: begin
				__main___storak17 <= convert_sync_array_muxed1;
			end
			5'd18: begin
				__main___storak18 <= convert_sync_array_muxed1;
			end
			5'd19: begin
				__main___storak19 <= convert_sync_array_muxed1;
			end
			5'd20: begin
				__main___storak20 <= convert_sync_array_muxed1;
			end
			5'd21: begin
				__main___storak21 <= convert_sync_array_muxed1;
			end
			5'd22: begin
				__main___storak22 <= convert_sync_array_muxed1;
			end
			5'd23: begin
				__main___storak23 <= convert_sync_array_muxed1;
			end
			5'd24: begin
				__main___storak24 <= convert_sync_array_muxed1;
			end
			5'd25: begin
				__main___storak25 <= convert_sync_array_muxed1;
			end
			5'd26: begin
				__main___storak26 <= convert_sync_array_muxed1;
			end
			5'd27: begin
				__main___storak27 <= convert_sync_array_muxed1;
			end
			5'd28: begin
				__main___storak28 <= convert_sync_array_muxed1;
			end
			5'd29: begin
				__main___storak29 <= convert_sync_array_muxed1;
			end
			5'd30: begin
				__main___storak30 <= convert_sync_array_muxed1;
			end
			default: begin
				__main___storak31 <= convert_sync_array_muxed1;
			end
		endcase
	end
	if (convert_t_next_value_ce) begin
		convert_sync_array_muxed2 = convert_t_next_value;
		case (ADR_i)
			1'd0: begin
				__main___storak0 <= convert_sync_array_muxed2;
			end
			1'd1: begin
				__main___storak1 <= convert_sync_array_muxed2;
			end
			2'd2: begin
				__main___storak2 <= convert_sync_array_muxed2;
			end
			2'd3: begin
				__main___storak3 <= convert_sync_array_muxed2;
			end
			3'd4: begin
				__main___storak4 <= convert_sync_array_muxed2;
			end
			3'd5: begin
				__main___storak5 <= convert_sync_array_muxed2;
			end
			3'd6: begin
				__main___storak6 <= convert_sync_array_muxed2;
			end
			3'd7: begin
				__main___storak7 <= convert_sync_array_muxed2;
			end
			4'd8: begin
				__main___storak8 <= convert_sync_array_muxed2;
			end
			4'd9: begin
				__main___storak9 <= convert_sync_array_muxed2;
			end
			4'd10: begin
				__main___storak10 <= convert_sync_array_muxed2;
			end
			4'd11: begin
				__main___storak11 <= convert_sync_array_muxed2;
			end
			4'd12: begin
				__main___storak12 <= convert_sync_array_muxed2;
			end
			4'd13: begin
				__main___storak13 <= convert_sync_array_muxed2;
			end
			4'd14: begin
				__main___storak14 <= convert_sync_array_muxed2;
			end
			4'd15: begin
				__main___storak15 <= convert_sync_array_muxed2;
			end
			5'd16: begin
				__main___storak16 <= convert_sync_array_muxed2;
			end
			5'd17: begin
				__main___storak17 <= convert_sync_array_muxed2;
			end
			5'd18: begin
				__main___storak18 <= convert_sync_array_muxed2;
			end
			5'd19: begin
				__main___storak19 <= convert_sync_array_muxed2;
			end
			5'd20: begin
				__main___storak20 <= convert_sync_array_muxed2;
			end
			5'd21: begin
				__main___storak21 <= convert_sync_array_muxed2;
			end
			5'd22: begin
				__main___storak22 <= convert_sync_array_muxed2;
			end
			5'd23: begin
				__main___storak23 <= convert_sync_array_muxed2;
			end
			5'd24: begin
				__main___storak24 <= convert_sync_array_muxed2;
			end
			5'd25: begin
				__main___storak25 <= convert_sync_array_muxed2;
			end
			5'd26: begin
				__main___storak26 <= convert_sync_array_muxed2;
			end
			5'd27: begin
				__main___storak27 <= convert_sync_array_muxed2;
			end
			5'd28: begin
				__main___storak28 <= convert_sync_array_muxed2;
			end
			5'd29: begin
				__main___storak29 <= convert_sync_array_muxed2;
			end
			5'd30: begin
				__main___storak30 <= convert_sync_array_muxed2;
			end
			default: begin
				__main___storak31 <= convert_sync_array_muxed2;
			end
		endcase
	end
	if (convert_f_next_value_ce) begin
		convert_sync_array_muxed3 = convert_f_next_value;
		case (ADR_i)
			1'd0: begin
				__main___storav0 <= convert_sync_array_muxed3;
			end
			1'd1: begin
				__main___storav1 <= convert_sync_array_muxed3;
			end
			2'd2: begin
				__main___storav2 <= convert_sync_array_muxed3;
			end
			2'd3: begin
				__main___storav3 <= convert_sync_array_muxed3;
			end
			3'd4: begin
				__main___storav4 <= convert_sync_array_muxed3;
			end
			3'd5: begin
				__main___storav5 <= convert_sync_array_muxed3;
			end
			3'd6: begin
				__main___storav6 <= convert_sync_array_muxed3;
			end
			3'd7: begin
				__main___storav7 <= convert_sync_array_muxed3;
			end
			4'd8: begin
				__main___storav8 <= convert_sync_array_muxed3;
			end
			4'd9: begin
				__main___storav9 <= convert_sync_array_muxed3;
			end
			4'd10: begin
				__main___storav10 <= convert_sync_array_muxed3;
			end
			4'd11: begin
				__main___storav11 <= convert_sync_array_muxed3;
			end
			4'd12: begin
				__main___storav12 <= convert_sync_array_muxed3;
			end
			4'd13: begin
				__main___storav13 <= convert_sync_array_muxed3;
			end
			4'd14: begin
				__main___storav14 <= convert_sync_array_muxed3;
			end
			4'd15: begin
				__main___storav15 <= convert_sync_array_muxed3;
			end
			5'd16: begin
				__main___storav16 <= convert_sync_array_muxed3;
			end
			5'd17: begin
				__main___storav17 <= convert_sync_array_muxed3;
			end
			5'd18: begin
				__main___storav18 <= convert_sync_array_muxed3;
			end
			5'd19: begin
				__main___storav19 <= convert_sync_array_muxed3;
			end
			5'd20: begin
				__main___storav20 <= convert_sync_array_muxed3;
			end
			5'd21: begin
				__main___storav21 <= convert_sync_array_muxed3;
			end
			5'd22: begin
				__main___storav22 <= convert_sync_array_muxed3;
			end
			5'd23: begin
				__main___storav23 <= convert_sync_array_muxed3;
			end
			5'd24: begin
				__main___storav24 <= convert_sync_array_muxed3;
			end
			5'd25: begin
				__main___storav25 <= convert_sync_array_muxed3;
			end
			5'd26: begin
				__main___storav26 <= convert_sync_array_muxed3;
			end
			5'd27: begin
				__main___storav27 <= convert_sync_array_muxed3;
			end
			5'd28: begin
				__main___storav28 <= convert_sync_array_muxed3;
			end
			5'd29: begin
				__main___storav29 <= convert_sync_array_muxed3;
			end
			5'd30: begin
				__main___storav30 <= convert_sync_array_muxed3;
			end
			default: begin
				__main___storav31 <= convert_sync_array_muxed3;
			end
		endcase
	end
	if (sys_rst_1) begin
		DUP_o <= 1'd0;
		STALL_o <= 1'd0;
		ACK_o <= 1'd0;
		DAT_o <= 16'd0;
		__main___storak0 <= 16'd0;
		__main___storak1 <= 16'd0;
		__main___storak2 <= 16'd0;
		__main___storak3 <= 16'd0;
		__main___storak4 <= 16'd0;
		__main___storak5 <= 16'd0;
		__main___storak6 <= 16'd0;
		__main___storak7 <= 16'd0;
		__main___storak8 <= 16'd0;
		__main___storak9 <= 16'd0;
		__main___storak10 <= 16'd0;
		__main___storak11 <= 16'd0;
		__main___storak12 <= 16'd0;
		__main___storak13 <= 16'd0;
		__main___storak14 <= 16'd0;
		__main___storak15 <= 16'd0;
		__main___storak16 <= 16'd0;
		__main___storak17 <= 16'd0;
		__main___storak18 <= 16'd0;
		__main___storak19 <= 16'd0;
		__main___storak20 <= 16'd0;
		__main___storak21 <= 16'd0;
		__main___storak22 <= 16'd0;
		__main___storak23 <= 16'd0;
		__main___storak24 <= 16'd0;
		__main___storak25 <= 16'd0;
		__main___storak26 <= 16'd0;
		__main___storak27 <= 16'd0;
		__main___storak28 <= 16'd0;
		__main___storak29 <= 16'd0;
		__main___storak30 <= 16'd0;
		__main___storak31 <= 16'd0;
		__main___storav0 <= 16'd0;
		__main___storav1 <= 16'd0;
		__main___storav2 <= 16'd0;
		__main___storav3 <= 16'd0;
		__main___storav4 <= 16'd0;
		__main___storav5 <= 16'd0;
		__main___storav6 <= 16'd0;
		__main___storav7 <= 16'd0;
		__main___storav8 <= 16'd0;
		__main___storav9 <= 16'd0;
		__main___storav10 <= 16'd0;
		__main___storav11 <= 16'd0;
		__main___storav12 <= 16'd0;
		__main___storav13 <= 16'd0;
		__main___storav14 <= 16'd0;
		__main___storav15 <= 16'd0;
		__main___storav16 <= 16'd0;
		__main___storav17 <= 16'd0;
		__main___storav18 <= 16'd0;
		__main___storav19 <= 16'd0;
		__main___storav20 <= 16'd0;
		__main___storav21 <= 16'd0;
		__main___storav22 <= 16'd0;
		__main___storav23 <= 16'd0;
		__main___storav24 <= 16'd0;
		__main___storav25 <= 16'd0;
		__main___storav26 <= 16'd0;
		__main___storav27 <= 16'd0;
		__main___storav28 <= 16'd0;
		__main___storav29 <= 16'd0;
		__main___storav30 <= 16'd0;
		__main___storav31 <= 16'd0;
		__main___empty_location <= 16'd1;
		convert_state <= 2'd3;
	end
end

endmodule


