VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_keyvalue
  CLASS BLOCK ;
  FOREIGN wrapped_keyvalue ;
  ORIGIN 0.000 0.000 ;
  SIZE 240.000 BY 240.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 236.000 9.570 240.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 219.000 240.000 219.600 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 236.000 12.330 240.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 236.000 88.690 240.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 236.000 98.810 240.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 236.000 223.930 240.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 216.280 240.000 216.880 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 236.000 127.330 240.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 236.000 17.850 240.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 27.240 240.000 27.840 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 170.040 240.000 170.640 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 236.000 71.210 240.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 236.000 142.050 240.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 204.040 240.000 204.640 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 61.240 240.000 61.840 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 236.000 65.690 240.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 236.000 22.450 240.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 236.000 180.690 240.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 236.000 157.690 240.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 236.000 62.930 240.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 233.960 240.000 234.560 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 236.000 208.290 240.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 236.000 190.810 240.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 178.200 240.000 178.800 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 106.120 240.000 106.720 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 236.000 52.810 240.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 54.440 240.000 55.040 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 236.000 116.290 240.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 236.000 91.450 240.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 129.240 240.000 129.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 144.200 240.000 144.800 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 236.000 94.210 240.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 236.000 205.530 240.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 148.280 240.000 148.880 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 50.360 240.000 50.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 236.000 114.450 240.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 236.000 121.810 240.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 118.360 240.000 118.960 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 236.000 73.050 240.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 125.160 240.000 125.760 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 238.040 240.000 238.640 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 236.000 119.050 240.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 174.120 240.000 174.720 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 236.000 192.650 240.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 236.000 234.050 240.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 236.000 78.570 240.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 42.200 240.000 42.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 236.000 167.810 240.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 236.000 235.890 240.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 46.280 240.000 46.880 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 236.000 42.690 240.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 236.000 19.690 240.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 84.360 240.000 84.960 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 236.000 139.290 240.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 236.000 175.170 240.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 197.240 240.000 197.840 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 236.000 144.810 240.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 236.000 162.290 240.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 133.320 240.000 133.920 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 31.320 240.000 31.920 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 236.000 84.090 240.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 236.000 27.970 240.000 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 236.000 40.850 240.000 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 163.240 240.000 163.840 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 236.000 228.530 240.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 236.000 96.050 240.000 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 236.000 75.810 240.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 69.400 240.000 70.000 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 227.160 240.000 227.760 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 236.000 2.210 240.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 114.280 240.000 114.880 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 236.000 129.170 240.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 236.000 131.930 240.000 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 9.560 240.000 10.160 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 12.280 240.000 12.880 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 236.000 30.730 240.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 236.000 198.170 240.000 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 236.000 101.570 240.000 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 140.120 240.000 140.720 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 185.000 240.000 185.600 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 236.000 124.570 240.000 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 236.000 35.330 240.000 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 236.000 68.450 240.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 121.080 240.000 121.680 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 137.400 240.000 138.000 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 236.000 215.650 240.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 91.160 240.000 91.760 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 236.000 15.090 240.000 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 236.000 188.050 240.000 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 155.080 240.000 155.680 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 236.000 147.570 240.000 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 24.520 240.000 25.120 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 236.000 177.930 240.000 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 65.320 240.000 65.920 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 236.000 238.650 240.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 35.400 240.000 36.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 193.160 240.000 193.760 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 236.000 218.410 240.000 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 236.000 154.930 240.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 236.000 7.730 240.000 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 236.000 48.210 240.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 236.000 159.530 240.000 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 212.200 240.000 212.800 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 236.000 85.930 240.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 236.000 50.970 240.000 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 236.000 165.050 240.000 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 228.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 228.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 236.000 134.690 240.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 5.480 240.000 6.080 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 236.000 221.170 240.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 236.000 182.530 240.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 236.000 58.330 240.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 236.000 55.570 240.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 110.200 240.000 110.800 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 95.240 240.000 95.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 76.200 240.000 76.800 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 1.400 240.000 2.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 236.000 211.050 240.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 208.120 240.000 208.720 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 236.000 108.930 240.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 236.000 149.410 240.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 80.280 240.000 80.880 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 182.280 240.000 182.880 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 236.000 231.290 240.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 39.480 240.000 40.080 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 236.000 137.450 240.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 236.000 32.570 240.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 236.000 45.450 240.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 236.000 38.090 240.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 73.480 240.000 74.080 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 236.000 200.930 240.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 231.240 240.000 231.840 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 236.000 81.330 240.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 223.080 240.000 223.680 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 152.360 240.000 152.960 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 236.000 225.770 240.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 236.000 111.690 240.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 103.400 240.000 104.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 16.360 240.000 16.960 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 57.160 240.000 57.760 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 236.000 212.890 240.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 189.080 240.000 189.680 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 99.320 240.000 99.920 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 199.960 240.000 200.560 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 236.000 202.770 240.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 236.000 195.410 240.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 236.000 104.330 240.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 236.000 152.170 240.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 236.000 106.170 240.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 236.000 185.290 240.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 20.440 240.000 21.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 167.320 240.000 167.920 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 159.160 240.000 159.760 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 236.000 172.410 240.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 236.000 170.570 240.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 236.000 25.210 240.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 236.000 61.090 240.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 236.000 4.970 240.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 236.000 88.440 240.000 89.040 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 236.295 238.255 ;
      LAYER met1 ;
        RECT 0.070 10.240 236.355 238.300 ;
      LAYER met2 ;
        RECT 0.100 235.720 1.650 238.525 ;
        RECT 2.490 235.720 4.410 238.525 ;
        RECT 5.250 235.720 7.170 238.525 ;
        RECT 8.010 235.720 9.010 238.525 ;
        RECT 9.850 235.720 11.770 238.525 ;
        RECT 12.610 235.720 14.530 238.525 ;
        RECT 15.370 235.720 17.290 238.525 ;
        RECT 18.130 235.720 19.130 238.525 ;
        RECT 19.970 235.720 21.890 238.525 ;
        RECT 22.730 235.720 24.650 238.525 ;
        RECT 25.490 235.720 27.410 238.525 ;
        RECT 28.250 235.720 30.170 238.525 ;
        RECT 31.010 235.720 32.010 238.525 ;
        RECT 32.850 235.720 34.770 238.525 ;
        RECT 35.610 235.720 37.530 238.525 ;
        RECT 38.370 235.720 40.290 238.525 ;
        RECT 41.130 235.720 42.130 238.525 ;
        RECT 42.970 235.720 44.890 238.525 ;
        RECT 45.730 235.720 47.650 238.525 ;
        RECT 48.490 235.720 50.410 238.525 ;
        RECT 51.250 235.720 52.250 238.525 ;
        RECT 53.090 235.720 55.010 238.525 ;
        RECT 55.850 235.720 57.770 238.525 ;
        RECT 58.610 235.720 60.530 238.525 ;
        RECT 61.370 235.720 62.370 238.525 ;
        RECT 63.210 235.720 65.130 238.525 ;
        RECT 65.970 235.720 67.890 238.525 ;
        RECT 68.730 235.720 70.650 238.525 ;
        RECT 71.490 235.720 72.490 238.525 ;
        RECT 73.330 235.720 75.250 238.525 ;
        RECT 76.090 235.720 78.010 238.525 ;
        RECT 78.850 235.720 80.770 238.525 ;
        RECT 81.610 235.720 83.530 238.525 ;
        RECT 84.370 235.720 85.370 238.525 ;
        RECT 86.210 235.720 88.130 238.525 ;
        RECT 88.970 235.720 90.890 238.525 ;
        RECT 91.730 235.720 93.650 238.525 ;
        RECT 94.490 235.720 95.490 238.525 ;
        RECT 96.330 235.720 98.250 238.525 ;
        RECT 99.090 235.720 101.010 238.525 ;
        RECT 101.850 235.720 103.770 238.525 ;
        RECT 104.610 235.720 105.610 238.525 ;
        RECT 106.450 235.720 108.370 238.525 ;
        RECT 109.210 235.720 111.130 238.525 ;
        RECT 111.970 235.720 113.890 238.525 ;
        RECT 114.730 235.720 115.730 238.525 ;
        RECT 116.570 235.720 118.490 238.525 ;
        RECT 119.330 235.720 121.250 238.525 ;
        RECT 122.090 235.720 124.010 238.525 ;
        RECT 124.850 235.720 126.770 238.525 ;
        RECT 127.610 235.720 128.610 238.525 ;
        RECT 129.450 235.720 131.370 238.525 ;
        RECT 132.210 235.720 134.130 238.525 ;
        RECT 134.970 235.720 136.890 238.525 ;
        RECT 137.730 235.720 138.730 238.525 ;
        RECT 139.570 235.720 141.490 238.525 ;
        RECT 142.330 235.720 144.250 238.525 ;
        RECT 145.090 235.720 147.010 238.525 ;
        RECT 147.850 235.720 148.850 238.525 ;
        RECT 149.690 235.720 151.610 238.525 ;
        RECT 152.450 235.720 154.370 238.525 ;
        RECT 155.210 235.720 157.130 238.525 ;
        RECT 157.970 235.720 158.970 238.525 ;
        RECT 159.810 235.720 161.730 238.525 ;
        RECT 162.570 235.720 164.490 238.525 ;
        RECT 165.330 235.720 167.250 238.525 ;
        RECT 168.090 235.720 170.010 238.525 ;
        RECT 170.850 235.720 171.850 238.525 ;
        RECT 172.690 235.720 174.610 238.525 ;
        RECT 175.450 235.720 177.370 238.525 ;
        RECT 178.210 235.720 180.130 238.525 ;
        RECT 180.970 235.720 181.970 238.525 ;
        RECT 182.810 235.720 184.730 238.525 ;
        RECT 185.570 235.720 187.490 238.525 ;
        RECT 188.330 235.720 190.250 238.525 ;
        RECT 191.090 235.720 192.090 238.525 ;
        RECT 192.930 235.720 194.850 238.525 ;
        RECT 195.690 235.720 197.610 238.525 ;
        RECT 198.450 235.720 200.370 238.525 ;
        RECT 201.210 235.720 202.210 238.525 ;
        RECT 203.050 235.720 204.970 238.525 ;
        RECT 205.810 235.720 207.730 238.525 ;
        RECT 208.570 235.720 210.490 238.525 ;
        RECT 211.330 235.720 212.330 238.525 ;
        RECT 213.170 235.720 215.090 238.525 ;
        RECT 215.930 235.720 217.850 238.525 ;
        RECT 218.690 235.720 220.610 238.525 ;
        RECT 221.450 235.720 223.370 238.525 ;
        RECT 224.210 235.720 225.210 238.525 ;
        RECT 226.050 235.720 227.970 238.525 ;
        RECT 228.810 235.720 230.730 238.525 ;
        RECT 231.570 235.720 233.490 238.525 ;
        RECT 234.330 235.720 235.330 238.525 ;
        RECT 0.100 4.280 235.880 235.720 ;
        RECT 0.650 2.875 1.650 4.280 ;
        RECT 2.490 2.875 4.410 4.280 ;
        RECT 5.250 2.875 7.170 4.280 ;
        RECT 8.010 2.875 9.930 4.280 ;
        RECT 10.770 2.875 11.770 4.280 ;
        RECT 12.610 2.875 14.530 4.280 ;
        RECT 15.370 2.875 17.290 4.280 ;
        RECT 18.130 2.875 20.050 4.280 ;
        RECT 20.890 2.875 21.890 4.280 ;
        RECT 22.730 2.875 24.650 4.280 ;
        RECT 25.490 2.875 27.410 4.280 ;
        RECT 28.250 2.875 30.170 4.280 ;
        RECT 31.010 2.875 32.010 4.280 ;
        RECT 32.850 2.875 34.770 4.280 ;
        RECT 35.610 2.875 37.530 4.280 ;
        RECT 38.370 2.875 40.290 4.280 ;
        RECT 41.130 2.875 42.130 4.280 ;
        RECT 42.970 2.875 44.890 4.280 ;
        RECT 45.730 2.875 47.650 4.280 ;
        RECT 48.490 2.875 50.410 4.280 ;
        RECT 51.250 2.875 53.170 4.280 ;
        RECT 54.010 2.875 55.010 4.280 ;
        RECT 55.850 2.875 57.770 4.280 ;
        RECT 58.610 2.875 60.530 4.280 ;
        RECT 61.370 2.875 63.290 4.280 ;
        RECT 64.130 2.875 65.130 4.280 ;
        RECT 65.970 2.875 67.890 4.280 ;
        RECT 68.730 2.875 70.650 4.280 ;
        RECT 71.490 2.875 73.410 4.280 ;
        RECT 74.250 2.875 75.250 4.280 ;
        RECT 76.090 2.875 78.010 4.280 ;
        RECT 78.850 2.875 80.770 4.280 ;
        RECT 81.610 2.875 83.530 4.280 ;
        RECT 84.370 2.875 85.370 4.280 ;
        RECT 86.210 2.875 88.130 4.280 ;
        RECT 88.970 2.875 90.890 4.280 ;
        RECT 91.730 2.875 93.650 4.280 ;
        RECT 94.490 2.875 96.410 4.280 ;
        RECT 97.250 2.875 98.250 4.280 ;
        RECT 99.090 2.875 101.010 4.280 ;
        RECT 101.850 2.875 103.770 4.280 ;
        RECT 104.610 2.875 106.530 4.280 ;
        RECT 107.370 2.875 108.370 4.280 ;
        RECT 109.210 2.875 111.130 4.280 ;
        RECT 111.970 2.875 113.890 4.280 ;
        RECT 114.730 2.875 116.650 4.280 ;
        RECT 117.490 2.875 118.490 4.280 ;
        RECT 119.330 2.875 121.250 4.280 ;
        RECT 122.090 2.875 124.010 4.280 ;
        RECT 124.850 2.875 126.770 4.280 ;
        RECT 127.610 2.875 128.610 4.280 ;
        RECT 129.450 2.875 131.370 4.280 ;
        RECT 132.210 2.875 134.130 4.280 ;
        RECT 134.970 2.875 136.890 4.280 ;
        RECT 137.730 2.875 138.730 4.280 ;
        RECT 139.570 2.875 141.490 4.280 ;
        RECT 142.330 2.875 144.250 4.280 ;
        RECT 145.090 2.875 147.010 4.280 ;
        RECT 147.850 2.875 149.770 4.280 ;
        RECT 150.610 2.875 151.610 4.280 ;
        RECT 152.450 2.875 154.370 4.280 ;
        RECT 155.210 2.875 157.130 4.280 ;
        RECT 157.970 2.875 159.890 4.280 ;
        RECT 160.730 2.875 161.730 4.280 ;
        RECT 162.570 2.875 164.490 4.280 ;
        RECT 165.330 2.875 167.250 4.280 ;
        RECT 168.090 2.875 170.010 4.280 ;
        RECT 170.850 2.875 171.850 4.280 ;
        RECT 172.690 2.875 174.610 4.280 ;
        RECT 175.450 2.875 177.370 4.280 ;
        RECT 178.210 2.875 180.130 4.280 ;
        RECT 180.970 2.875 181.970 4.280 ;
        RECT 182.810 2.875 184.730 4.280 ;
        RECT 185.570 2.875 187.490 4.280 ;
        RECT 188.330 2.875 190.250 4.280 ;
        RECT 191.090 2.875 193.010 4.280 ;
        RECT 193.850 2.875 194.850 4.280 ;
        RECT 195.690 2.875 197.610 4.280 ;
        RECT 198.450 2.875 200.370 4.280 ;
        RECT 201.210 2.875 203.130 4.280 ;
        RECT 203.970 2.875 204.970 4.280 ;
        RECT 205.810 2.875 207.730 4.280 ;
        RECT 208.570 2.875 210.490 4.280 ;
        RECT 211.330 2.875 213.250 4.280 ;
        RECT 214.090 2.875 215.090 4.280 ;
        RECT 215.930 2.875 217.850 4.280 ;
        RECT 218.690 2.875 220.610 4.280 ;
        RECT 221.450 2.875 223.370 4.280 ;
        RECT 224.210 2.875 225.210 4.280 ;
        RECT 226.050 2.875 227.970 4.280 ;
        RECT 228.810 2.875 230.730 4.280 ;
        RECT 231.570 2.875 233.490 4.280 ;
        RECT 234.330 2.875 235.330 4.280 ;
      LAYER met3 ;
        RECT 4.000 237.680 235.600 238.505 ;
        RECT 4.400 237.640 235.600 237.680 ;
        RECT 4.400 236.280 236.000 237.640 ;
        RECT 4.000 234.960 236.000 236.280 ;
        RECT 4.000 233.600 235.600 234.960 ;
        RECT 4.400 233.560 235.600 233.600 ;
        RECT 4.400 232.240 236.000 233.560 ;
        RECT 4.400 232.200 235.600 232.240 ;
        RECT 4.000 230.840 235.600 232.200 ;
        RECT 4.000 229.520 236.000 230.840 ;
        RECT 4.400 228.160 236.000 229.520 ;
        RECT 4.400 228.120 235.600 228.160 ;
        RECT 4.000 226.760 235.600 228.120 ;
        RECT 4.000 225.440 236.000 226.760 ;
        RECT 4.400 224.080 236.000 225.440 ;
        RECT 4.400 224.040 235.600 224.080 ;
        RECT 4.000 222.720 235.600 224.040 ;
        RECT 4.400 222.680 235.600 222.720 ;
        RECT 4.400 221.320 236.000 222.680 ;
        RECT 4.000 220.000 236.000 221.320 ;
        RECT 4.000 218.640 235.600 220.000 ;
        RECT 4.400 218.600 235.600 218.640 ;
        RECT 4.400 217.280 236.000 218.600 ;
        RECT 4.400 217.240 235.600 217.280 ;
        RECT 4.000 215.880 235.600 217.240 ;
        RECT 4.000 214.560 236.000 215.880 ;
        RECT 4.400 213.200 236.000 214.560 ;
        RECT 4.400 213.160 235.600 213.200 ;
        RECT 4.000 211.800 235.600 213.160 ;
        RECT 4.000 210.480 236.000 211.800 ;
        RECT 4.400 209.120 236.000 210.480 ;
        RECT 4.400 209.080 235.600 209.120 ;
        RECT 4.000 207.720 235.600 209.080 ;
        RECT 4.000 206.400 236.000 207.720 ;
        RECT 4.400 205.040 236.000 206.400 ;
        RECT 4.400 205.000 235.600 205.040 ;
        RECT 4.000 203.680 235.600 205.000 ;
        RECT 4.400 203.640 235.600 203.680 ;
        RECT 4.400 202.280 236.000 203.640 ;
        RECT 4.000 200.960 236.000 202.280 ;
        RECT 4.000 199.600 235.600 200.960 ;
        RECT 4.400 199.560 235.600 199.600 ;
        RECT 4.400 198.240 236.000 199.560 ;
        RECT 4.400 198.200 235.600 198.240 ;
        RECT 4.000 196.840 235.600 198.200 ;
        RECT 4.000 195.520 236.000 196.840 ;
        RECT 4.400 194.160 236.000 195.520 ;
        RECT 4.400 194.120 235.600 194.160 ;
        RECT 4.000 192.760 235.600 194.120 ;
        RECT 4.000 191.440 236.000 192.760 ;
        RECT 4.400 190.080 236.000 191.440 ;
        RECT 4.400 190.040 235.600 190.080 ;
        RECT 4.000 188.720 235.600 190.040 ;
        RECT 4.400 188.680 235.600 188.720 ;
        RECT 4.400 187.320 236.000 188.680 ;
        RECT 4.000 186.000 236.000 187.320 ;
        RECT 4.000 184.640 235.600 186.000 ;
        RECT 4.400 184.600 235.600 184.640 ;
        RECT 4.400 183.280 236.000 184.600 ;
        RECT 4.400 183.240 235.600 183.280 ;
        RECT 4.000 181.880 235.600 183.240 ;
        RECT 4.000 180.560 236.000 181.880 ;
        RECT 4.400 179.200 236.000 180.560 ;
        RECT 4.400 179.160 235.600 179.200 ;
        RECT 4.000 177.800 235.600 179.160 ;
        RECT 4.000 176.480 236.000 177.800 ;
        RECT 4.400 175.120 236.000 176.480 ;
        RECT 4.400 175.080 235.600 175.120 ;
        RECT 4.000 173.760 235.600 175.080 ;
        RECT 4.400 173.720 235.600 173.760 ;
        RECT 4.400 172.360 236.000 173.720 ;
        RECT 4.000 171.040 236.000 172.360 ;
        RECT 4.000 169.680 235.600 171.040 ;
        RECT 4.400 169.640 235.600 169.680 ;
        RECT 4.400 168.320 236.000 169.640 ;
        RECT 4.400 168.280 235.600 168.320 ;
        RECT 4.000 166.920 235.600 168.280 ;
        RECT 4.000 165.600 236.000 166.920 ;
        RECT 4.400 164.240 236.000 165.600 ;
        RECT 4.400 164.200 235.600 164.240 ;
        RECT 4.000 162.840 235.600 164.200 ;
        RECT 4.000 161.520 236.000 162.840 ;
        RECT 4.400 160.160 236.000 161.520 ;
        RECT 4.400 160.120 235.600 160.160 ;
        RECT 4.000 158.800 235.600 160.120 ;
        RECT 4.400 158.760 235.600 158.800 ;
        RECT 4.400 157.400 236.000 158.760 ;
        RECT 4.000 156.080 236.000 157.400 ;
        RECT 4.000 154.720 235.600 156.080 ;
        RECT 4.400 154.680 235.600 154.720 ;
        RECT 4.400 153.360 236.000 154.680 ;
        RECT 4.400 153.320 235.600 153.360 ;
        RECT 4.000 151.960 235.600 153.320 ;
        RECT 4.000 150.640 236.000 151.960 ;
        RECT 4.400 149.280 236.000 150.640 ;
        RECT 4.400 149.240 235.600 149.280 ;
        RECT 4.000 147.880 235.600 149.240 ;
        RECT 4.000 146.560 236.000 147.880 ;
        RECT 4.400 145.200 236.000 146.560 ;
        RECT 4.400 145.160 235.600 145.200 ;
        RECT 4.000 143.840 235.600 145.160 ;
        RECT 4.400 143.800 235.600 143.840 ;
        RECT 4.400 142.440 236.000 143.800 ;
        RECT 4.000 141.120 236.000 142.440 ;
        RECT 4.000 139.760 235.600 141.120 ;
        RECT 4.400 139.720 235.600 139.760 ;
        RECT 4.400 138.400 236.000 139.720 ;
        RECT 4.400 138.360 235.600 138.400 ;
        RECT 4.000 137.000 235.600 138.360 ;
        RECT 4.000 135.680 236.000 137.000 ;
        RECT 4.400 134.320 236.000 135.680 ;
        RECT 4.400 134.280 235.600 134.320 ;
        RECT 4.000 132.920 235.600 134.280 ;
        RECT 4.000 131.600 236.000 132.920 ;
        RECT 4.400 130.240 236.000 131.600 ;
        RECT 4.400 130.200 235.600 130.240 ;
        RECT 4.000 128.840 235.600 130.200 ;
        RECT 4.000 127.520 236.000 128.840 ;
        RECT 4.400 126.160 236.000 127.520 ;
        RECT 4.400 126.120 235.600 126.160 ;
        RECT 4.000 124.800 235.600 126.120 ;
        RECT 4.400 124.760 235.600 124.800 ;
        RECT 4.400 123.400 236.000 124.760 ;
        RECT 4.000 122.080 236.000 123.400 ;
        RECT 4.000 120.720 235.600 122.080 ;
        RECT 4.400 120.680 235.600 120.720 ;
        RECT 4.400 119.360 236.000 120.680 ;
        RECT 4.400 119.320 235.600 119.360 ;
        RECT 4.000 117.960 235.600 119.320 ;
        RECT 4.000 116.640 236.000 117.960 ;
        RECT 4.400 115.280 236.000 116.640 ;
        RECT 4.400 115.240 235.600 115.280 ;
        RECT 4.000 113.880 235.600 115.240 ;
        RECT 4.000 112.560 236.000 113.880 ;
        RECT 4.400 111.200 236.000 112.560 ;
        RECT 4.400 111.160 235.600 111.200 ;
        RECT 4.000 109.840 235.600 111.160 ;
        RECT 4.400 109.800 235.600 109.840 ;
        RECT 4.400 108.440 236.000 109.800 ;
        RECT 4.000 107.120 236.000 108.440 ;
        RECT 4.000 105.760 235.600 107.120 ;
        RECT 4.400 105.720 235.600 105.760 ;
        RECT 4.400 104.400 236.000 105.720 ;
        RECT 4.400 104.360 235.600 104.400 ;
        RECT 4.000 103.000 235.600 104.360 ;
        RECT 4.000 101.680 236.000 103.000 ;
        RECT 4.400 100.320 236.000 101.680 ;
        RECT 4.400 100.280 235.600 100.320 ;
        RECT 4.000 98.920 235.600 100.280 ;
        RECT 4.000 97.600 236.000 98.920 ;
        RECT 4.400 96.240 236.000 97.600 ;
        RECT 4.400 96.200 235.600 96.240 ;
        RECT 4.000 94.880 235.600 96.200 ;
        RECT 4.400 94.840 235.600 94.880 ;
        RECT 4.400 93.480 236.000 94.840 ;
        RECT 4.000 92.160 236.000 93.480 ;
        RECT 4.000 90.800 235.600 92.160 ;
        RECT 4.400 90.760 235.600 90.800 ;
        RECT 4.400 89.440 236.000 90.760 ;
        RECT 4.400 89.400 235.600 89.440 ;
        RECT 4.000 88.040 235.600 89.400 ;
        RECT 4.000 86.720 236.000 88.040 ;
        RECT 4.400 85.360 236.000 86.720 ;
        RECT 4.400 85.320 235.600 85.360 ;
        RECT 4.000 83.960 235.600 85.320 ;
        RECT 4.000 82.640 236.000 83.960 ;
        RECT 4.400 81.280 236.000 82.640 ;
        RECT 4.400 81.240 235.600 81.280 ;
        RECT 4.000 79.920 235.600 81.240 ;
        RECT 4.400 79.880 235.600 79.920 ;
        RECT 4.400 78.520 236.000 79.880 ;
        RECT 4.000 77.200 236.000 78.520 ;
        RECT 4.000 75.840 235.600 77.200 ;
        RECT 4.400 75.800 235.600 75.840 ;
        RECT 4.400 74.480 236.000 75.800 ;
        RECT 4.400 74.440 235.600 74.480 ;
        RECT 4.000 73.080 235.600 74.440 ;
        RECT 4.000 71.760 236.000 73.080 ;
        RECT 4.400 70.400 236.000 71.760 ;
        RECT 4.400 70.360 235.600 70.400 ;
        RECT 4.000 69.000 235.600 70.360 ;
        RECT 4.000 67.680 236.000 69.000 ;
        RECT 4.400 66.320 236.000 67.680 ;
        RECT 4.400 66.280 235.600 66.320 ;
        RECT 4.000 64.920 235.600 66.280 ;
        RECT 4.000 63.600 236.000 64.920 ;
        RECT 4.400 62.240 236.000 63.600 ;
        RECT 4.400 62.200 235.600 62.240 ;
        RECT 4.000 60.880 235.600 62.200 ;
        RECT 4.400 60.840 235.600 60.880 ;
        RECT 4.400 59.480 236.000 60.840 ;
        RECT 4.000 58.160 236.000 59.480 ;
        RECT 4.000 56.800 235.600 58.160 ;
        RECT 4.400 56.760 235.600 56.800 ;
        RECT 4.400 55.440 236.000 56.760 ;
        RECT 4.400 55.400 235.600 55.440 ;
        RECT 4.000 54.040 235.600 55.400 ;
        RECT 4.000 52.720 236.000 54.040 ;
        RECT 4.400 51.360 236.000 52.720 ;
        RECT 4.400 51.320 235.600 51.360 ;
        RECT 4.000 49.960 235.600 51.320 ;
        RECT 4.000 48.640 236.000 49.960 ;
        RECT 4.400 47.280 236.000 48.640 ;
        RECT 4.400 47.240 235.600 47.280 ;
        RECT 4.000 45.920 235.600 47.240 ;
        RECT 4.400 45.880 235.600 45.920 ;
        RECT 4.400 44.520 236.000 45.880 ;
        RECT 4.000 43.200 236.000 44.520 ;
        RECT 4.000 41.840 235.600 43.200 ;
        RECT 4.400 41.800 235.600 41.840 ;
        RECT 4.400 40.480 236.000 41.800 ;
        RECT 4.400 40.440 235.600 40.480 ;
        RECT 4.000 39.080 235.600 40.440 ;
        RECT 4.000 37.760 236.000 39.080 ;
        RECT 4.400 36.400 236.000 37.760 ;
        RECT 4.400 36.360 235.600 36.400 ;
        RECT 4.000 35.000 235.600 36.360 ;
        RECT 4.000 33.680 236.000 35.000 ;
        RECT 4.400 32.320 236.000 33.680 ;
        RECT 4.400 32.280 235.600 32.320 ;
        RECT 4.000 30.960 235.600 32.280 ;
        RECT 4.400 30.920 235.600 30.960 ;
        RECT 4.400 29.560 236.000 30.920 ;
        RECT 4.000 28.240 236.000 29.560 ;
        RECT 4.000 26.880 235.600 28.240 ;
        RECT 4.400 26.840 235.600 26.880 ;
        RECT 4.400 25.520 236.000 26.840 ;
        RECT 4.400 25.480 235.600 25.520 ;
        RECT 4.000 24.120 235.600 25.480 ;
        RECT 4.000 22.800 236.000 24.120 ;
        RECT 4.400 21.440 236.000 22.800 ;
        RECT 4.400 21.400 235.600 21.440 ;
        RECT 4.000 20.040 235.600 21.400 ;
        RECT 4.000 18.720 236.000 20.040 ;
        RECT 4.400 17.360 236.000 18.720 ;
        RECT 4.400 17.320 235.600 17.360 ;
        RECT 4.000 16.000 235.600 17.320 ;
        RECT 4.400 15.960 235.600 16.000 ;
        RECT 4.400 14.600 236.000 15.960 ;
        RECT 4.000 13.280 236.000 14.600 ;
        RECT 4.000 11.920 235.600 13.280 ;
        RECT 4.400 11.880 235.600 11.920 ;
        RECT 4.400 10.560 236.000 11.880 ;
        RECT 4.400 10.520 235.600 10.560 ;
        RECT 4.000 9.160 235.600 10.520 ;
        RECT 4.000 7.840 236.000 9.160 ;
        RECT 4.400 6.480 236.000 7.840 ;
        RECT 4.400 6.440 235.600 6.480 ;
        RECT 4.000 5.080 235.600 6.440 ;
        RECT 4.000 3.760 236.000 5.080 ;
        RECT 4.400 2.895 236.000 3.760 ;
      LAYER met4 ;
        RECT 100.575 96.735 100.905 114.065 ;
  END
END wrapped_keyvalue
END LIBRARY

