/* Machine-generated using Migen */
module keyvalue_3(
	input sys_rst,
	input [3:0] SEL_i,
	input ADR_IS_KEY_i,
	input DAT_IS_KEY_i,
	input [63:0] ADR_i,
	input [63:0] DAT_i,
	input WE_i,
	input STB_i,
	input CYC_i,
	input DUP_o,
	output reg STALL_o,
	output reg ACK_o,
	output reg [63:0] DAT_o,
	output [63:0] LA_o,
	input sys_clk,
	input sys_rst_1
);

reg [63:0] __main___storak0 = 64'd0;
reg [63:0] __main___storak1 = 64'd0;
reg [63:0] __main___storak2 = 64'd0;
reg [63:0] __main___storak3 = 64'd0;
reg [63:0] __main___storak4 = 64'd0;
reg [63:0] __main___storak5 = 64'd0;
reg [63:0] __main___storak6 = 64'd0;
reg [63:0] __main___storak7 = 64'd0;
reg [63:0] __main___storak8 = 64'd0;
reg [63:0] __main___storak9 = 64'd0;
reg [63:0] __main___storak10 = 64'd0;
reg [63:0] __main___storak11 = 64'd0;
reg [63:0] __main___storak12 = 64'd0;
reg [63:0] __main___storak13 = 64'd0;
reg [63:0] __main___storak14 = 64'd0;
reg [63:0] __main___storak15 = 64'd0;
reg [63:0] __main___storak16 = 64'd0;
reg [63:0] __main___storak17 = 64'd0;
reg [63:0] __main___storak18 = 64'd0;
reg [63:0] __main___storak19 = 64'd0;
reg [63:0] __main___storak20 = 64'd0;
reg [63:0] __main___storak21 = 64'd0;
reg [63:0] __main___storak22 = 64'd0;
reg [63:0] __main___storak23 = 64'd0;
reg [63:0] __main___storak24 = 64'd0;
reg [63:0] __main___storak25 = 64'd0;
reg [63:0] __main___storak26 = 64'd0;
reg [63:0] __main___storak27 = 64'd0;
reg [63:0] __main___storak28 = 64'd0;
reg [63:0] __main___storak29 = 64'd0;
reg [63:0] __main___storak30 = 64'd0;
reg [63:0] __main___storak31 = 64'd0;
reg [63:0] __main___storak32 = 64'd0;
reg [63:0] __main___storak33 = 64'd0;
reg [63:0] __main___storak34 = 64'd0;
reg [63:0] __main___storak35 = 64'd0;
reg [63:0] __main___storak36 = 64'd0;
reg [63:0] __main___storak37 = 64'd0;
reg [63:0] __main___storak38 = 64'd0;
reg [63:0] __main___storak39 = 64'd0;
reg [63:0] __main___storak40 = 64'd0;
reg [63:0] __main___storak41 = 64'd0;
reg [63:0] __main___storak42 = 64'd0;
reg [63:0] __main___storak43 = 64'd0;
reg [63:0] __main___storak44 = 64'd0;
reg [63:0] __main___storak45 = 64'd0;
reg [63:0] __main___storak46 = 64'd0;
reg [63:0] __main___storak47 = 64'd0;
reg [63:0] __main___storak48 = 64'd0;
reg [63:0] __main___storak49 = 64'd0;
reg [63:0] __main___storak50 = 64'd0;
reg [63:0] __main___storak51 = 64'd0;
reg [63:0] __main___storak52 = 64'd0;
reg [63:0] __main___storak53 = 64'd0;
reg [63:0] __main___storak54 = 64'd0;
reg [63:0] __main___storak55 = 64'd0;
reg [63:0] __main___storak56 = 64'd0;
reg [63:0] __main___storak57 = 64'd0;
reg [63:0] __main___storak58 = 64'd0;
reg [63:0] __main___storak59 = 64'd0;
reg [63:0] __main___storak60 = 64'd0;
reg [63:0] __main___storak61 = 64'd0;
reg [63:0] __main___storak62 = 64'd0;
reg [63:0] __main___storak63 = 64'd0;
reg [63:0] __main___storak64 = 64'd0;
reg [63:0] __main___storak65 = 64'd0;
reg [63:0] __main___storak66 = 64'd0;
reg [63:0] __main___storak67 = 64'd0;
reg [63:0] __main___storak68 = 64'd0;
reg [63:0] __main___storak69 = 64'd0;
reg [63:0] __main___storak70 = 64'd0;
reg [63:0] __main___storak71 = 64'd0;
reg [63:0] __main___storak72 = 64'd0;
reg [63:0] __main___storak73 = 64'd0;
reg [63:0] __main___storak74 = 64'd0;
reg [63:0] __main___storak75 = 64'd0;
reg [63:0] __main___storak76 = 64'd0;
reg [63:0] __main___storak77 = 64'd0;
reg [63:0] __main___storak78 = 64'd0;
reg [63:0] __main___storak79 = 64'd0;
reg [63:0] __main___storak80 = 64'd0;
reg [63:0] __main___storak81 = 64'd0;
reg [63:0] __main___storak82 = 64'd0;
reg [63:0] __main___storak83 = 64'd0;
reg [63:0] __main___storak84 = 64'd0;
reg [63:0] __main___storak85 = 64'd0;
reg [63:0] __main___storak86 = 64'd0;
reg [63:0] __main___storak87 = 64'd0;
reg [63:0] __main___storak88 = 64'd0;
reg [63:0] __main___storak89 = 64'd0;
reg [63:0] __main___storak90 = 64'd0;
reg [63:0] __main___storak91 = 64'd0;
reg [63:0] __main___storak92 = 64'd0;
reg [63:0] __main___storak93 = 64'd0;
reg [63:0] __main___storak94 = 64'd0;
reg [63:0] __main___storak95 = 64'd0;
reg [63:0] __main___storak96 = 64'd0;
reg [63:0] __main___storak97 = 64'd0;
reg [63:0] __main___storak98 = 64'd0;
reg [63:0] __main___storak99 = 64'd0;
reg [63:0] __main___storak100 = 64'd0;
reg [63:0] __main___storak101 = 64'd0;
reg [63:0] __main___storak102 = 64'd0;
reg [63:0] __main___storak103 = 64'd0;
reg [63:0] __main___storak104 = 64'd0;
reg [63:0] __main___storak105 = 64'd0;
reg [63:0] __main___storak106 = 64'd0;
reg [63:0] __main___storak107 = 64'd0;
reg [63:0] __main___storak108 = 64'd0;
reg [63:0] __main___storak109 = 64'd0;
reg [63:0] __main___storak110 = 64'd0;
reg [63:0] __main___storak111 = 64'd0;
reg [63:0] __main___storak112 = 64'd0;
reg [63:0] __main___storak113 = 64'd0;
reg [63:0] __main___storak114 = 64'd0;
reg [63:0] __main___storak115 = 64'd0;
reg [63:0] __main___storak116 = 64'd0;
reg [63:0] __main___storak117 = 64'd0;
reg [63:0] __main___storak118 = 64'd0;
reg [63:0] __main___storak119 = 64'd0;
reg [63:0] __main___storak120 = 64'd0;
reg [63:0] __main___storak121 = 64'd0;
reg [63:0] __main___storak122 = 64'd0;
reg [63:0] __main___storak123 = 64'd0;
reg [63:0] __main___storak124 = 64'd0;
reg [63:0] __main___storak125 = 64'd0;
reg [63:0] __main___storak126 = 64'd0;
reg [63:0] __main___storak127 = 64'd0;
reg [63:0] __main___storav0 = 64'd0;
reg [63:0] __main___storav1 = 64'd0;
reg [63:0] __main___storav2 = 64'd0;
reg [63:0] __main___storav3 = 64'd0;
reg [63:0] __main___storav4 = 64'd0;
reg [63:0] __main___storav5 = 64'd0;
reg [63:0] __main___storav6 = 64'd0;
reg [63:0] __main___storav7 = 64'd0;
reg [63:0] __main___storav8 = 64'd0;
reg [63:0] __main___storav9 = 64'd0;
reg [63:0] __main___storav10 = 64'd0;
reg [63:0] __main___storav11 = 64'd0;
reg [63:0] __main___storav12 = 64'd0;
reg [63:0] __main___storav13 = 64'd0;
reg [63:0] __main___storav14 = 64'd0;
reg [63:0] __main___storav15 = 64'd0;
reg [63:0] __main___storav16 = 64'd0;
reg [63:0] __main___storav17 = 64'd0;
reg [63:0] __main___storav18 = 64'd0;
reg [63:0] __main___storav19 = 64'd0;
reg [63:0] __main___storav20 = 64'd0;
reg [63:0] __main___storav21 = 64'd0;
reg [63:0] __main___storav22 = 64'd0;
reg [63:0] __main___storav23 = 64'd0;
reg [63:0] __main___storav24 = 64'd0;
reg [63:0] __main___storav25 = 64'd0;
reg [63:0] __main___storav26 = 64'd0;
reg [63:0] __main___storav27 = 64'd0;
reg [63:0] __main___storav28 = 64'd0;
reg [63:0] __main___storav29 = 64'd0;
reg [63:0] __main___storav30 = 64'd0;
reg [63:0] __main___storav31 = 64'd0;
reg [63:0] __main___storav32 = 64'd0;
reg [63:0] __main___storav33 = 64'd0;
reg [63:0] __main___storav34 = 64'd0;
reg [63:0] __main___storav35 = 64'd0;
reg [63:0] __main___storav36 = 64'd0;
reg [63:0] __main___storav37 = 64'd0;
reg [63:0] __main___storav38 = 64'd0;
reg [63:0] __main___storav39 = 64'd0;
reg [63:0] __main___storav40 = 64'd0;
reg [63:0] __main___storav41 = 64'd0;
reg [63:0] __main___storav42 = 64'd0;
reg [63:0] __main___storav43 = 64'd0;
reg [63:0] __main___storav44 = 64'd0;
reg [63:0] __main___storav45 = 64'd0;
reg [63:0] __main___storav46 = 64'd0;
reg [63:0] __main___storav47 = 64'd0;
reg [63:0] __main___storav48 = 64'd0;
reg [63:0] __main___storav49 = 64'd0;
reg [63:0] __main___storav50 = 64'd0;
reg [63:0] __main___storav51 = 64'd0;
reg [63:0] __main___storav52 = 64'd0;
reg [63:0] __main___storav53 = 64'd0;
reg [63:0] __main___storav54 = 64'd0;
reg [63:0] __main___storav55 = 64'd0;
reg [63:0] __main___storav56 = 64'd0;
reg [63:0] __main___storav57 = 64'd0;
reg [63:0] __main___storav58 = 64'd0;
reg [63:0] __main___storav59 = 64'd0;
reg [63:0] __main___storav60 = 64'd0;
reg [63:0] __main___storav61 = 64'd0;
reg [63:0] __main___storav62 = 64'd0;
reg [63:0] __main___storav63 = 64'd0;
reg [63:0] __main___storav64 = 64'd0;
reg [63:0] __main___storav65 = 64'd0;
reg [63:0] __main___storav66 = 64'd0;
reg [63:0] __main___storav67 = 64'd0;
reg [63:0] __main___storav68 = 64'd0;
reg [63:0] __main___storav69 = 64'd0;
reg [63:0] __main___storav70 = 64'd0;
reg [63:0] __main___storav71 = 64'd0;
reg [63:0] __main___storav72 = 64'd0;
reg [63:0] __main___storav73 = 64'd0;
reg [63:0] __main___storav74 = 64'd0;
reg [63:0] __main___storav75 = 64'd0;
reg [63:0] __main___storav76 = 64'd0;
reg [63:0] __main___storav77 = 64'd0;
reg [63:0] __main___storav78 = 64'd0;
reg [63:0] __main___storav79 = 64'd0;
reg [63:0] __main___storav80 = 64'd0;
reg [63:0] __main___storav81 = 64'd0;
reg [63:0] __main___storav82 = 64'd0;
reg [63:0] __main___storav83 = 64'd0;
reg [63:0] __main___storav84 = 64'd0;
reg [63:0] __main___storav85 = 64'd0;
reg [63:0] __main___storav86 = 64'd0;
reg [63:0] __main___storav87 = 64'd0;
reg [63:0] __main___storav88 = 64'd0;
reg [63:0] __main___storav89 = 64'd0;
reg [63:0] __main___storav90 = 64'd0;
reg [63:0] __main___storav91 = 64'd0;
reg [63:0] __main___storav92 = 64'd0;
reg [63:0] __main___storav93 = 64'd0;
reg [63:0] __main___storav94 = 64'd0;
reg [63:0] __main___storav95 = 64'd0;
reg [63:0] __main___storav96 = 64'd0;
reg [63:0] __main___storav97 = 64'd0;
reg [63:0] __main___storav98 = 64'd0;
reg [63:0] __main___storav99 = 64'd0;
reg [63:0] __main___storav100 = 64'd0;
reg [63:0] __main___storav101 = 64'd0;
reg [63:0] __main___storav102 = 64'd0;
reg [63:0] __main___storav103 = 64'd0;
reg [63:0] __main___storav104 = 64'd0;
reg [63:0] __main___storav105 = 64'd0;
reg [63:0] __main___storav106 = 64'd0;
reg [63:0] __main___storav107 = 64'd0;
reg [63:0] __main___storav108 = 64'd0;
reg [63:0] __main___storav109 = 64'd0;
reg [63:0] __main___storav110 = 64'd0;
reg [63:0] __main___storav111 = 64'd0;
reg [63:0] __main___storav112 = 64'd0;
reg [63:0] __main___storav113 = 64'd0;
reg [63:0] __main___storav114 = 64'd0;
reg [63:0] __main___storav115 = 64'd0;
reg [63:0] __main___storav116 = 64'd0;
reg [63:0] __main___storav117 = 64'd0;
reg [63:0] __main___storav118 = 64'd0;
reg [63:0] __main___storav119 = 64'd0;
reg [63:0] __main___storav120 = 64'd0;
reg [63:0] __main___storav121 = 64'd0;
reg [63:0] __main___storav122 = 64'd0;
reg [63:0] __main___storav123 = 64'd0;
reg [63:0] __main___storav124 = 64'd0;
reg [63:0] __main___storav125 = 64'd0;
reg [63:0] __main___storav126 = 64'd0;
reg [63:0] __main___storav127 = 64'd0;
reg [63:0] __main___empty_location = 64'd0;
reg [1:0] convert_state = 2'd3;
reg [1:0] convert_next_state;
reg __main___STALL_o_next_value0;
reg __main___STALL_o_next_value_ce0;
reg [63:0] __main___empty_location_t_next_value;
reg __main___empty_location_t_next_value_ce;
reg __main___ACK_o_f_next_value;
reg __main___ACK_o_f_next_value_ce;
reg [63:0] __main___DAT_o_next_value1;
reg __main___DAT_o_next_value_ce1;
reg [63:0] convert_next_value0;
reg convert_next_value_ce0;
reg [63:0] convert_next_value1;
reg convert_next_value_ce1;
reg [63:0] convert_t_next_value;
reg convert_t_next_value_ce;
reg [63:0] convert_f_next_value;
reg convert_f_next_value_ce;
reg [63:0] convert_comb_array_muxed;
reg [63:0] convert_sync_array_muxed0 = 64'd0;
reg [63:0] convert_sync_array_muxed1 = 64'd0;
reg [63:0] convert_sync_array_muxed2 = 64'd0;
reg [63:0] convert_sync_array_muxed3 = 64'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign LA_o = DAT_o;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	convert_next_state <= 2'd0;
	__main___STALL_o_next_value0 <= 1'd0;
	__main___STALL_o_next_value_ce0 <= 1'd0;
	__main___empty_location_t_next_value <= 64'd0;
	__main___empty_location_t_next_value_ce <= 1'd0;
	__main___ACK_o_f_next_value <= 1'd0;
	__main___ACK_o_f_next_value_ce <= 1'd0;
	__main___DAT_o_next_value1 <= 64'd0;
	__main___DAT_o_next_value_ce1 <= 1'd0;
	convert_next_value0 <= 64'd0;
	convert_next_value_ce0 <= 1'd0;
	convert_next_value1 <= 64'd0;
	convert_next_value_ce1 <= 1'd0;
	convert_t_next_value <= 64'd0;
	convert_t_next_value_ce <= 1'd0;
	convert_f_next_value <= 64'd0;
	convert_f_next_value_ce <= 1'd0;
	convert_next_state <= convert_state;
	case (convert_state)
		1'd0: begin
			__main___STALL_o_next_value0 <= 1'd0;
			__main___STALL_o_next_value_ce0 <= 1'd1;
			if ((((STB_i == 1'd1) & (WE_i == 1'd0)) & (ACK_o == 1'd0))) begin
				convert_next_state <= 1'd1;
			end else begin
				if ((((STB_i == 1'd1) & (WE_i == 1'd1)) & (ACK_o == 1'd0))) begin
					convert_next_state <= 2'd2;
					if ((ADR_i == 64'd0)) begin
						__main___empty_location_t_next_value <= (__main___empty_location + 1'd1);
						__main___empty_location_t_next_value_ce <= 1'd1;
					end
				end else begin
					__main___ACK_o_f_next_value <= 1'd0;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
		end
		1'd1: begin
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak1 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav1;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak2 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav2;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak3 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav3;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak4 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav4;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak5 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav5;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak6 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav6;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak7 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav7;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak8 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav8;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak9 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav9;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak10 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav10;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak11 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav11;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak12 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav12;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak13 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav13;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak14 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav14;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak15 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav15;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak16 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav16;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak17 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav17;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak18 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav18;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak19 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav19;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak20 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav20;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak21 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav21;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak22 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav22;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak23 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav23;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak24 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav24;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak25 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav25;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak26 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav26;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak27 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav27;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak28 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav28;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak29 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav29;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak30 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav30;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak31 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav31;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak32 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav32;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak33 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav33;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak34 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav34;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak35 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav35;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak36 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav36;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak37 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav37;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak38 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav38;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak39 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav39;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak40 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav40;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak41 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav41;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak42 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav42;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak43 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav43;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak44 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav44;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak45 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav45;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak46 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav46;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak47 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav47;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak48 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav48;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak49 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav49;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak50 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav50;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak51 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav51;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak52 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav52;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak53 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav53;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak54 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav54;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak55 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav55;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak56 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav56;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak57 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav57;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak58 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav58;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak59 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav59;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak60 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav60;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak61 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav61;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak62 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav62;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak63 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav63;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak64 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav64;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak65 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav65;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak66 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav66;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak67 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav67;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak68 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav68;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak69 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav69;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak70 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav70;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak71 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav71;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak72 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav72;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak73 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav73;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak74 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav74;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak75 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav75;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak76 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav76;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak77 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav77;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak78 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav78;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak79 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav79;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak80 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav80;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak81 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav81;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak82 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav82;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak83 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav83;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak84 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav84;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak85 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav85;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak86 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav86;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak87 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav87;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak88 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav88;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak89 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav89;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak90 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav90;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak91 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav91;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak92 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav92;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak93 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav93;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak94 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav94;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak95 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav95;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak96 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav96;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak97 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav97;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak98 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav98;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak99 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav99;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak100 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav100;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak101 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav101;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak102 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav102;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak103 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav103;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak104 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav104;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak105 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav105;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak106 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav106;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak107 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav107;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak108 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav108;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak109 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav109;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak110 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav110;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak111 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav111;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak112 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav112;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak113 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav113;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak114 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav114;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak115 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav115;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak116 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav116;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak117 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav117;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak118 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav118;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak119 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav119;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak120 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav120;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak121 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav121;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak122 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav122;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak123 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav123;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak124 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav124;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak125 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav125;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak126 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav126;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd1)) begin
				if ((__main___storak127 == ADR_i)) begin
					__main___DAT_o_next_value1 <= __main___storav127;
					__main___DAT_o_next_value_ce1 <= 1'd1;
					__main___ACK_o_f_next_value <= 1'd1;
					__main___ACK_o_f_next_value_ce <= 1'd1;
					convert_next_state <= 1'd0;
				end
			end
			if ((ADR_IS_KEY_i == 1'd0)) begin
				__main___DAT_o_next_value1 <= convert_comb_array_muxed;
				__main___DAT_o_next_value_ce1 <= 1'd1;
				__main___ACK_o_f_next_value <= 1'd1;
				__main___ACK_o_f_next_value_ce <= 1'd1;
				convert_next_state <= 1'd0;
			end
			if ((sys_rst == 1'd1)) begin
				convert_next_state <= 2'd3;
			end
		end
		2'd2: begin
			if (ADR_IS_KEY_i) begin
				convert_next_value0 <= DAT_i;
				convert_next_value_ce0 <= 1'd1;
				convert_next_value1 <= ADR_i;
				convert_next_value_ce1 <= 1'd1;
				__main___DAT_o_next_value1 <= __main___empty_location;
				__main___DAT_o_next_value_ce1 <= 1'd1;
			end else begin
				if (DAT_IS_KEY_i) begin
					convert_t_next_value <= DAT_i;
					convert_t_next_value_ce <= 1'd1;
					__main___DAT_o_next_value1 <= ADR_i;
					__main___DAT_o_next_value_ce1 <= 1'd1;
				end else begin
					convert_f_next_value <= DAT_i;
					convert_f_next_value_ce <= 1'd1;
					__main___DAT_o_next_value1 <= ADR_i;
					__main___DAT_o_next_value_ce1 <= 1'd1;
				end
			end
			__main___ACK_o_f_next_value <= 1'd1;
			__main___ACK_o_f_next_value_ce <= 1'd1;
			convert_next_state <= 1'd0;
			if ((sys_rst == 1'd1)) begin
				convert_next_state <= 2'd3;
			end else begin
				convert_next_state <= 1'd0;
			end
		end
		default: begin
			convert_next_state <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	convert_comb_array_muxed <= 64'd0;
	case (ADR_i)
		1'd0: begin
			convert_comb_array_muxed <= __main___storav0;
		end
		1'd1: begin
			convert_comb_array_muxed <= __main___storav1;
		end
		2'd2: begin
			convert_comb_array_muxed <= __main___storav2;
		end
		2'd3: begin
			convert_comb_array_muxed <= __main___storav3;
		end
		3'd4: begin
			convert_comb_array_muxed <= __main___storav4;
		end
		3'd5: begin
			convert_comb_array_muxed <= __main___storav5;
		end
		3'd6: begin
			convert_comb_array_muxed <= __main___storav6;
		end
		3'd7: begin
			convert_comb_array_muxed <= __main___storav7;
		end
		4'd8: begin
			convert_comb_array_muxed <= __main___storav8;
		end
		4'd9: begin
			convert_comb_array_muxed <= __main___storav9;
		end
		4'd10: begin
			convert_comb_array_muxed <= __main___storav10;
		end
		4'd11: begin
			convert_comb_array_muxed <= __main___storav11;
		end
		4'd12: begin
			convert_comb_array_muxed <= __main___storav12;
		end
		4'd13: begin
			convert_comb_array_muxed <= __main___storav13;
		end
		4'd14: begin
			convert_comb_array_muxed <= __main___storav14;
		end
		4'd15: begin
			convert_comb_array_muxed <= __main___storav15;
		end
		5'd16: begin
			convert_comb_array_muxed <= __main___storav16;
		end
		5'd17: begin
			convert_comb_array_muxed <= __main___storav17;
		end
		5'd18: begin
			convert_comb_array_muxed <= __main___storav18;
		end
		5'd19: begin
			convert_comb_array_muxed <= __main___storav19;
		end
		5'd20: begin
			convert_comb_array_muxed <= __main___storav20;
		end
		5'd21: begin
			convert_comb_array_muxed <= __main___storav21;
		end
		5'd22: begin
			convert_comb_array_muxed <= __main___storav22;
		end
		5'd23: begin
			convert_comb_array_muxed <= __main___storav23;
		end
		5'd24: begin
			convert_comb_array_muxed <= __main___storav24;
		end
		5'd25: begin
			convert_comb_array_muxed <= __main___storav25;
		end
		5'd26: begin
			convert_comb_array_muxed <= __main___storav26;
		end
		5'd27: begin
			convert_comb_array_muxed <= __main___storav27;
		end
		5'd28: begin
			convert_comb_array_muxed <= __main___storav28;
		end
		5'd29: begin
			convert_comb_array_muxed <= __main___storav29;
		end
		5'd30: begin
			convert_comb_array_muxed <= __main___storav30;
		end
		5'd31: begin
			convert_comb_array_muxed <= __main___storav31;
		end
		6'd32: begin
			convert_comb_array_muxed <= __main___storav32;
		end
		6'd33: begin
			convert_comb_array_muxed <= __main___storav33;
		end
		6'd34: begin
			convert_comb_array_muxed <= __main___storav34;
		end
		6'd35: begin
			convert_comb_array_muxed <= __main___storav35;
		end
		6'd36: begin
			convert_comb_array_muxed <= __main___storav36;
		end
		6'd37: begin
			convert_comb_array_muxed <= __main___storav37;
		end
		6'd38: begin
			convert_comb_array_muxed <= __main___storav38;
		end
		6'd39: begin
			convert_comb_array_muxed <= __main___storav39;
		end
		6'd40: begin
			convert_comb_array_muxed <= __main___storav40;
		end
		6'd41: begin
			convert_comb_array_muxed <= __main___storav41;
		end
		6'd42: begin
			convert_comb_array_muxed <= __main___storav42;
		end
		6'd43: begin
			convert_comb_array_muxed <= __main___storav43;
		end
		6'd44: begin
			convert_comb_array_muxed <= __main___storav44;
		end
		6'd45: begin
			convert_comb_array_muxed <= __main___storav45;
		end
		6'd46: begin
			convert_comb_array_muxed <= __main___storav46;
		end
		6'd47: begin
			convert_comb_array_muxed <= __main___storav47;
		end
		6'd48: begin
			convert_comb_array_muxed <= __main___storav48;
		end
		6'd49: begin
			convert_comb_array_muxed <= __main___storav49;
		end
		6'd50: begin
			convert_comb_array_muxed <= __main___storav50;
		end
		6'd51: begin
			convert_comb_array_muxed <= __main___storav51;
		end
		6'd52: begin
			convert_comb_array_muxed <= __main___storav52;
		end
		6'd53: begin
			convert_comb_array_muxed <= __main___storav53;
		end
		6'd54: begin
			convert_comb_array_muxed <= __main___storav54;
		end
		6'd55: begin
			convert_comb_array_muxed <= __main___storav55;
		end
		6'd56: begin
			convert_comb_array_muxed <= __main___storav56;
		end
		6'd57: begin
			convert_comb_array_muxed <= __main___storav57;
		end
		6'd58: begin
			convert_comb_array_muxed <= __main___storav58;
		end
		6'd59: begin
			convert_comb_array_muxed <= __main___storav59;
		end
		6'd60: begin
			convert_comb_array_muxed <= __main___storav60;
		end
		6'd61: begin
			convert_comb_array_muxed <= __main___storav61;
		end
		6'd62: begin
			convert_comb_array_muxed <= __main___storav62;
		end
		6'd63: begin
			convert_comb_array_muxed <= __main___storav63;
		end
		7'd64: begin
			convert_comb_array_muxed <= __main___storav64;
		end
		7'd65: begin
			convert_comb_array_muxed <= __main___storav65;
		end
		7'd66: begin
			convert_comb_array_muxed <= __main___storav66;
		end
		7'd67: begin
			convert_comb_array_muxed <= __main___storav67;
		end
		7'd68: begin
			convert_comb_array_muxed <= __main___storav68;
		end
		7'd69: begin
			convert_comb_array_muxed <= __main___storav69;
		end
		7'd70: begin
			convert_comb_array_muxed <= __main___storav70;
		end
		7'd71: begin
			convert_comb_array_muxed <= __main___storav71;
		end
		7'd72: begin
			convert_comb_array_muxed <= __main___storav72;
		end
		7'd73: begin
			convert_comb_array_muxed <= __main___storav73;
		end
		7'd74: begin
			convert_comb_array_muxed <= __main___storav74;
		end
		7'd75: begin
			convert_comb_array_muxed <= __main___storav75;
		end
		7'd76: begin
			convert_comb_array_muxed <= __main___storav76;
		end
		7'd77: begin
			convert_comb_array_muxed <= __main___storav77;
		end
		7'd78: begin
			convert_comb_array_muxed <= __main___storav78;
		end
		7'd79: begin
			convert_comb_array_muxed <= __main___storav79;
		end
		7'd80: begin
			convert_comb_array_muxed <= __main___storav80;
		end
		7'd81: begin
			convert_comb_array_muxed <= __main___storav81;
		end
		7'd82: begin
			convert_comb_array_muxed <= __main___storav82;
		end
		7'd83: begin
			convert_comb_array_muxed <= __main___storav83;
		end
		7'd84: begin
			convert_comb_array_muxed <= __main___storav84;
		end
		7'd85: begin
			convert_comb_array_muxed <= __main___storav85;
		end
		7'd86: begin
			convert_comb_array_muxed <= __main___storav86;
		end
		7'd87: begin
			convert_comb_array_muxed <= __main___storav87;
		end
		7'd88: begin
			convert_comb_array_muxed <= __main___storav88;
		end
		7'd89: begin
			convert_comb_array_muxed <= __main___storav89;
		end
		7'd90: begin
			convert_comb_array_muxed <= __main___storav90;
		end
		7'd91: begin
			convert_comb_array_muxed <= __main___storav91;
		end
		7'd92: begin
			convert_comb_array_muxed <= __main___storav92;
		end
		7'd93: begin
			convert_comb_array_muxed <= __main___storav93;
		end
		7'd94: begin
			convert_comb_array_muxed <= __main___storav94;
		end
		7'd95: begin
			convert_comb_array_muxed <= __main___storav95;
		end
		7'd96: begin
			convert_comb_array_muxed <= __main___storav96;
		end
		7'd97: begin
			convert_comb_array_muxed <= __main___storav97;
		end
		7'd98: begin
			convert_comb_array_muxed <= __main___storav98;
		end
		7'd99: begin
			convert_comb_array_muxed <= __main___storav99;
		end
		7'd100: begin
			convert_comb_array_muxed <= __main___storav100;
		end
		7'd101: begin
			convert_comb_array_muxed <= __main___storav101;
		end
		7'd102: begin
			convert_comb_array_muxed <= __main___storav102;
		end
		7'd103: begin
			convert_comb_array_muxed <= __main___storav103;
		end
		7'd104: begin
			convert_comb_array_muxed <= __main___storav104;
		end
		7'd105: begin
			convert_comb_array_muxed <= __main___storav105;
		end
		7'd106: begin
			convert_comb_array_muxed <= __main___storav106;
		end
		7'd107: begin
			convert_comb_array_muxed <= __main___storav107;
		end
		7'd108: begin
			convert_comb_array_muxed <= __main___storav108;
		end
		7'd109: begin
			convert_comb_array_muxed <= __main___storav109;
		end
		7'd110: begin
			convert_comb_array_muxed <= __main___storav110;
		end
		7'd111: begin
			convert_comb_array_muxed <= __main___storav111;
		end
		7'd112: begin
			convert_comb_array_muxed <= __main___storav112;
		end
		7'd113: begin
			convert_comb_array_muxed <= __main___storav113;
		end
		7'd114: begin
			convert_comb_array_muxed <= __main___storav114;
		end
		7'd115: begin
			convert_comb_array_muxed <= __main___storav115;
		end
		7'd116: begin
			convert_comb_array_muxed <= __main___storav116;
		end
		7'd117: begin
			convert_comb_array_muxed <= __main___storav117;
		end
		7'd118: begin
			convert_comb_array_muxed <= __main___storav118;
		end
		7'd119: begin
			convert_comb_array_muxed <= __main___storav119;
		end
		7'd120: begin
			convert_comb_array_muxed <= __main___storav120;
		end
		7'd121: begin
			convert_comb_array_muxed <= __main___storav121;
		end
		7'd122: begin
			convert_comb_array_muxed <= __main___storav122;
		end
		7'd123: begin
			convert_comb_array_muxed <= __main___storav123;
		end
		7'd124: begin
			convert_comb_array_muxed <= __main___storav124;
		end
		7'd125: begin
			convert_comb_array_muxed <= __main___storav125;
		end
		7'd126: begin
			convert_comb_array_muxed <= __main___storav126;
		end
		default: begin
			convert_comb_array_muxed <= __main___storav127;
		end
	endcase
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

always @(posedge sys_clk) begin
	convert_state <= convert_next_state;
	if (__main___STALL_o_next_value_ce0) begin
		STALL_o <= __main___STALL_o_next_value0;
	end
	if (__main___empty_location_t_next_value_ce) begin
		__main___empty_location <= __main___empty_location_t_next_value;
	end
	if (__main___ACK_o_f_next_value_ce) begin
		ACK_o <= __main___ACK_o_f_next_value;
	end
	if (__main___DAT_o_next_value_ce1) begin
		DAT_o <= __main___DAT_o_next_value1;
	end
	if (convert_next_value_ce0) begin
		convert_sync_array_muxed0 = convert_next_value0;
		case (__main___empty_location)
			1'd0: begin
				__main___storav0 <= convert_sync_array_muxed0;
			end
			1'd1: begin
				__main___storav1 <= convert_sync_array_muxed0;
			end
			2'd2: begin
				__main___storav2 <= convert_sync_array_muxed0;
			end
			2'd3: begin
				__main___storav3 <= convert_sync_array_muxed0;
			end
			3'd4: begin
				__main___storav4 <= convert_sync_array_muxed0;
			end
			3'd5: begin
				__main___storav5 <= convert_sync_array_muxed0;
			end
			3'd6: begin
				__main___storav6 <= convert_sync_array_muxed0;
			end
			3'd7: begin
				__main___storav7 <= convert_sync_array_muxed0;
			end
			4'd8: begin
				__main___storav8 <= convert_sync_array_muxed0;
			end
			4'd9: begin
				__main___storav9 <= convert_sync_array_muxed0;
			end
			4'd10: begin
				__main___storav10 <= convert_sync_array_muxed0;
			end
			4'd11: begin
				__main___storav11 <= convert_sync_array_muxed0;
			end
			4'd12: begin
				__main___storav12 <= convert_sync_array_muxed0;
			end
			4'd13: begin
				__main___storav13 <= convert_sync_array_muxed0;
			end
			4'd14: begin
				__main___storav14 <= convert_sync_array_muxed0;
			end
			4'd15: begin
				__main___storav15 <= convert_sync_array_muxed0;
			end
			5'd16: begin
				__main___storav16 <= convert_sync_array_muxed0;
			end
			5'd17: begin
				__main___storav17 <= convert_sync_array_muxed0;
			end
			5'd18: begin
				__main___storav18 <= convert_sync_array_muxed0;
			end
			5'd19: begin
				__main___storav19 <= convert_sync_array_muxed0;
			end
			5'd20: begin
				__main___storav20 <= convert_sync_array_muxed0;
			end
			5'd21: begin
				__main___storav21 <= convert_sync_array_muxed0;
			end
			5'd22: begin
				__main___storav22 <= convert_sync_array_muxed0;
			end
			5'd23: begin
				__main___storav23 <= convert_sync_array_muxed0;
			end
			5'd24: begin
				__main___storav24 <= convert_sync_array_muxed0;
			end
			5'd25: begin
				__main___storav25 <= convert_sync_array_muxed0;
			end
			5'd26: begin
				__main___storav26 <= convert_sync_array_muxed0;
			end
			5'd27: begin
				__main___storav27 <= convert_sync_array_muxed0;
			end
			5'd28: begin
				__main___storav28 <= convert_sync_array_muxed0;
			end
			5'd29: begin
				__main___storav29 <= convert_sync_array_muxed0;
			end
			5'd30: begin
				__main___storav30 <= convert_sync_array_muxed0;
			end
			5'd31: begin
				__main___storav31 <= convert_sync_array_muxed0;
			end
			6'd32: begin
				__main___storav32 <= convert_sync_array_muxed0;
			end
			6'd33: begin
				__main___storav33 <= convert_sync_array_muxed0;
			end
			6'd34: begin
				__main___storav34 <= convert_sync_array_muxed0;
			end
			6'd35: begin
				__main___storav35 <= convert_sync_array_muxed0;
			end
			6'd36: begin
				__main___storav36 <= convert_sync_array_muxed0;
			end
			6'd37: begin
				__main___storav37 <= convert_sync_array_muxed0;
			end
			6'd38: begin
				__main___storav38 <= convert_sync_array_muxed0;
			end
			6'd39: begin
				__main___storav39 <= convert_sync_array_muxed0;
			end
			6'd40: begin
				__main___storav40 <= convert_sync_array_muxed0;
			end
			6'd41: begin
				__main___storav41 <= convert_sync_array_muxed0;
			end
			6'd42: begin
				__main___storav42 <= convert_sync_array_muxed0;
			end
			6'd43: begin
				__main___storav43 <= convert_sync_array_muxed0;
			end
			6'd44: begin
				__main___storav44 <= convert_sync_array_muxed0;
			end
			6'd45: begin
				__main___storav45 <= convert_sync_array_muxed0;
			end
			6'd46: begin
				__main___storav46 <= convert_sync_array_muxed0;
			end
			6'd47: begin
				__main___storav47 <= convert_sync_array_muxed0;
			end
			6'd48: begin
				__main___storav48 <= convert_sync_array_muxed0;
			end
			6'd49: begin
				__main___storav49 <= convert_sync_array_muxed0;
			end
			6'd50: begin
				__main___storav50 <= convert_sync_array_muxed0;
			end
			6'd51: begin
				__main___storav51 <= convert_sync_array_muxed0;
			end
			6'd52: begin
				__main___storav52 <= convert_sync_array_muxed0;
			end
			6'd53: begin
				__main___storav53 <= convert_sync_array_muxed0;
			end
			6'd54: begin
				__main___storav54 <= convert_sync_array_muxed0;
			end
			6'd55: begin
				__main___storav55 <= convert_sync_array_muxed0;
			end
			6'd56: begin
				__main___storav56 <= convert_sync_array_muxed0;
			end
			6'd57: begin
				__main___storav57 <= convert_sync_array_muxed0;
			end
			6'd58: begin
				__main___storav58 <= convert_sync_array_muxed0;
			end
			6'd59: begin
				__main___storav59 <= convert_sync_array_muxed0;
			end
			6'd60: begin
				__main___storav60 <= convert_sync_array_muxed0;
			end
			6'd61: begin
				__main___storav61 <= convert_sync_array_muxed0;
			end
			6'd62: begin
				__main___storav62 <= convert_sync_array_muxed0;
			end
			6'd63: begin
				__main___storav63 <= convert_sync_array_muxed0;
			end
			7'd64: begin
				__main___storav64 <= convert_sync_array_muxed0;
			end
			7'd65: begin
				__main___storav65 <= convert_sync_array_muxed0;
			end
			7'd66: begin
				__main___storav66 <= convert_sync_array_muxed0;
			end
			7'd67: begin
				__main___storav67 <= convert_sync_array_muxed0;
			end
			7'd68: begin
				__main___storav68 <= convert_sync_array_muxed0;
			end
			7'd69: begin
				__main___storav69 <= convert_sync_array_muxed0;
			end
			7'd70: begin
				__main___storav70 <= convert_sync_array_muxed0;
			end
			7'd71: begin
				__main___storav71 <= convert_sync_array_muxed0;
			end
			7'd72: begin
				__main___storav72 <= convert_sync_array_muxed0;
			end
			7'd73: begin
				__main___storav73 <= convert_sync_array_muxed0;
			end
			7'd74: begin
				__main___storav74 <= convert_sync_array_muxed0;
			end
			7'd75: begin
				__main___storav75 <= convert_sync_array_muxed0;
			end
			7'd76: begin
				__main___storav76 <= convert_sync_array_muxed0;
			end
			7'd77: begin
				__main___storav77 <= convert_sync_array_muxed0;
			end
			7'd78: begin
				__main___storav78 <= convert_sync_array_muxed0;
			end
			7'd79: begin
				__main___storav79 <= convert_sync_array_muxed0;
			end
			7'd80: begin
				__main___storav80 <= convert_sync_array_muxed0;
			end
			7'd81: begin
				__main___storav81 <= convert_sync_array_muxed0;
			end
			7'd82: begin
				__main___storav82 <= convert_sync_array_muxed0;
			end
			7'd83: begin
				__main___storav83 <= convert_sync_array_muxed0;
			end
			7'd84: begin
				__main___storav84 <= convert_sync_array_muxed0;
			end
			7'd85: begin
				__main___storav85 <= convert_sync_array_muxed0;
			end
			7'd86: begin
				__main___storav86 <= convert_sync_array_muxed0;
			end
			7'd87: begin
				__main___storav87 <= convert_sync_array_muxed0;
			end
			7'd88: begin
				__main___storav88 <= convert_sync_array_muxed0;
			end
			7'd89: begin
				__main___storav89 <= convert_sync_array_muxed0;
			end
			7'd90: begin
				__main___storav90 <= convert_sync_array_muxed0;
			end
			7'd91: begin
				__main___storav91 <= convert_sync_array_muxed0;
			end
			7'd92: begin
				__main___storav92 <= convert_sync_array_muxed0;
			end
			7'd93: begin
				__main___storav93 <= convert_sync_array_muxed0;
			end
			7'd94: begin
				__main___storav94 <= convert_sync_array_muxed0;
			end
			7'd95: begin
				__main___storav95 <= convert_sync_array_muxed0;
			end
			7'd96: begin
				__main___storav96 <= convert_sync_array_muxed0;
			end
			7'd97: begin
				__main___storav97 <= convert_sync_array_muxed0;
			end
			7'd98: begin
				__main___storav98 <= convert_sync_array_muxed0;
			end
			7'd99: begin
				__main___storav99 <= convert_sync_array_muxed0;
			end
			7'd100: begin
				__main___storav100 <= convert_sync_array_muxed0;
			end
			7'd101: begin
				__main___storav101 <= convert_sync_array_muxed0;
			end
			7'd102: begin
				__main___storav102 <= convert_sync_array_muxed0;
			end
			7'd103: begin
				__main___storav103 <= convert_sync_array_muxed0;
			end
			7'd104: begin
				__main___storav104 <= convert_sync_array_muxed0;
			end
			7'd105: begin
				__main___storav105 <= convert_sync_array_muxed0;
			end
			7'd106: begin
				__main___storav106 <= convert_sync_array_muxed0;
			end
			7'd107: begin
				__main___storav107 <= convert_sync_array_muxed0;
			end
			7'd108: begin
				__main___storav108 <= convert_sync_array_muxed0;
			end
			7'd109: begin
				__main___storav109 <= convert_sync_array_muxed0;
			end
			7'd110: begin
				__main___storav110 <= convert_sync_array_muxed0;
			end
			7'd111: begin
				__main___storav111 <= convert_sync_array_muxed0;
			end
			7'd112: begin
				__main___storav112 <= convert_sync_array_muxed0;
			end
			7'd113: begin
				__main___storav113 <= convert_sync_array_muxed0;
			end
			7'd114: begin
				__main___storav114 <= convert_sync_array_muxed0;
			end
			7'd115: begin
				__main___storav115 <= convert_sync_array_muxed0;
			end
			7'd116: begin
				__main___storav116 <= convert_sync_array_muxed0;
			end
			7'd117: begin
				__main___storav117 <= convert_sync_array_muxed0;
			end
			7'd118: begin
				__main___storav118 <= convert_sync_array_muxed0;
			end
			7'd119: begin
				__main___storav119 <= convert_sync_array_muxed0;
			end
			7'd120: begin
				__main___storav120 <= convert_sync_array_muxed0;
			end
			7'd121: begin
				__main___storav121 <= convert_sync_array_muxed0;
			end
			7'd122: begin
				__main___storav122 <= convert_sync_array_muxed0;
			end
			7'd123: begin
				__main___storav123 <= convert_sync_array_muxed0;
			end
			7'd124: begin
				__main___storav124 <= convert_sync_array_muxed0;
			end
			7'd125: begin
				__main___storav125 <= convert_sync_array_muxed0;
			end
			7'd126: begin
				__main___storav126 <= convert_sync_array_muxed0;
			end
			default: begin
				__main___storav127 <= convert_sync_array_muxed0;
			end
		endcase
	end
	if (convert_next_value_ce1) begin
		convert_sync_array_muxed1 = convert_next_value1;
		case (__main___empty_location)
			1'd0: begin
				__main___storak0 <= convert_sync_array_muxed1;
			end
			1'd1: begin
				__main___storak1 <= convert_sync_array_muxed1;
			end
			2'd2: begin
				__main___storak2 <= convert_sync_array_muxed1;
			end
			2'd3: begin
				__main___storak3 <= convert_sync_array_muxed1;
			end
			3'd4: begin
				__main___storak4 <= convert_sync_array_muxed1;
			end
			3'd5: begin
				__main___storak5 <= convert_sync_array_muxed1;
			end
			3'd6: begin
				__main___storak6 <= convert_sync_array_muxed1;
			end
			3'd7: begin
				__main___storak7 <= convert_sync_array_muxed1;
			end
			4'd8: begin
				__main___storak8 <= convert_sync_array_muxed1;
			end
			4'd9: begin
				__main___storak9 <= convert_sync_array_muxed1;
			end
			4'd10: begin
				__main___storak10 <= convert_sync_array_muxed1;
			end
			4'd11: begin
				__main___storak11 <= convert_sync_array_muxed1;
			end
			4'd12: begin
				__main___storak12 <= convert_sync_array_muxed1;
			end
			4'd13: begin
				__main___storak13 <= convert_sync_array_muxed1;
			end
			4'd14: begin
				__main___storak14 <= convert_sync_array_muxed1;
			end
			4'd15: begin
				__main___storak15 <= convert_sync_array_muxed1;
			end
			5'd16: begin
				__main___storak16 <= convert_sync_array_muxed1;
			end
			5'd17: begin
				__main___storak17 <= convert_sync_array_muxed1;
			end
			5'd18: begin
				__main___storak18 <= convert_sync_array_muxed1;
			end
			5'd19: begin
				__main___storak19 <= convert_sync_array_muxed1;
			end
			5'd20: begin
				__main___storak20 <= convert_sync_array_muxed1;
			end
			5'd21: begin
				__main___storak21 <= convert_sync_array_muxed1;
			end
			5'd22: begin
				__main___storak22 <= convert_sync_array_muxed1;
			end
			5'd23: begin
				__main___storak23 <= convert_sync_array_muxed1;
			end
			5'd24: begin
				__main___storak24 <= convert_sync_array_muxed1;
			end
			5'd25: begin
				__main___storak25 <= convert_sync_array_muxed1;
			end
			5'd26: begin
				__main___storak26 <= convert_sync_array_muxed1;
			end
			5'd27: begin
				__main___storak27 <= convert_sync_array_muxed1;
			end
			5'd28: begin
				__main___storak28 <= convert_sync_array_muxed1;
			end
			5'd29: begin
				__main___storak29 <= convert_sync_array_muxed1;
			end
			5'd30: begin
				__main___storak30 <= convert_sync_array_muxed1;
			end
			5'd31: begin
				__main___storak31 <= convert_sync_array_muxed1;
			end
			6'd32: begin
				__main___storak32 <= convert_sync_array_muxed1;
			end
			6'd33: begin
				__main___storak33 <= convert_sync_array_muxed1;
			end
			6'd34: begin
				__main___storak34 <= convert_sync_array_muxed1;
			end
			6'd35: begin
				__main___storak35 <= convert_sync_array_muxed1;
			end
			6'd36: begin
				__main___storak36 <= convert_sync_array_muxed1;
			end
			6'd37: begin
				__main___storak37 <= convert_sync_array_muxed1;
			end
			6'd38: begin
				__main___storak38 <= convert_sync_array_muxed1;
			end
			6'd39: begin
				__main___storak39 <= convert_sync_array_muxed1;
			end
			6'd40: begin
				__main___storak40 <= convert_sync_array_muxed1;
			end
			6'd41: begin
				__main___storak41 <= convert_sync_array_muxed1;
			end
			6'd42: begin
				__main___storak42 <= convert_sync_array_muxed1;
			end
			6'd43: begin
				__main___storak43 <= convert_sync_array_muxed1;
			end
			6'd44: begin
				__main___storak44 <= convert_sync_array_muxed1;
			end
			6'd45: begin
				__main___storak45 <= convert_sync_array_muxed1;
			end
			6'd46: begin
				__main___storak46 <= convert_sync_array_muxed1;
			end
			6'd47: begin
				__main___storak47 <= convert_sync_array_muxed1;
			end
			6'd48: begin
				__main___storak48 <= convert_sync_array_muxed1;
			end
			6'd49: begin
				__main___storak49 <= convert_sync_array_muxed1;
			end
			6'd50: begin
				__main___storak50 <= convert_sync_array_muxed1;
			end
			6'd51: begin
				__main___storak51 <= convert_sync_array_muxed1;
			end
			6'd52: begin
				__main___storak52 <= convert_sync_array_muxed1;
			end
			6'd53: begin
				__main___storak53 <= convert_sync_array_muxed1;
			end
			6'd54: begin
				__main___storak54 <= convert_sync_array_muxed1;
			end
			6'd55: begin
				__main___storak55 <= convert_sync_array_muxed1;
			end
			6'd56: begin
				__main___storak56 <= convert_sync_array_muxed1;
			end
			6'd57: begin
				__main___storak57 <= convert_sync_array_muxed1;
			end
			6'd58: begin
				__main___storak58 <= convert_sync_array_muxed1;
			end
			6'd59: begin
				__main___storak59 <= convert_sync_array_muxed1;
			end
			6'd60: begin
				__main___storak60 <= convert_sync_array_muxed1;
			end
			6'd61: begin
				__main___storak61 <= convert_sync_array_muxed1;
			end
			6'd62: begin
				__main___storak62 <= convert_sync_array_muxed1;
			end
			6'd63: begin
				__main___storak63 <= convert_sync_array_muxed1;
			end
			7'd64: begin
				__main___storak64 <= convert_sync_array_muxed1;
			end
			7'd65: begin
				__main___storak65 <= convert_sync_array_muxed1;
			end
			7'd66: begin
				__main___storak66 <= convert_sync_array_muxed1;
			end
			7'd67: begin
				__main___storak67 <= convert_sync_array_muxed1;
			end
			7'd68: begin
				__main___storak68 <= convert_sync_array_muxed1;
			end
			7'd69: begin
				__main___storak69 <= convert_sync_array_muxed1;
			end
			7'd70: begin
				__main___storak70 <= convert_sync_array_muxed1;
			end
			7'd71: begin
				__main___storak71 <= convert_sync_array_muxed1;
			end
			7'd72: begin
				__main___storak72 <= convert_sync_array_muxed1;
			end
			7'd73: begin
				__main___storak73 <= convert_sync_array_muxed1;
			end
			7'd74: begin
				__main___storak74 <= convert_sync_array_muxed1;
			end
			7'd75: begin
				__main___storak75 <= convert_sync_array_muxed1;
			end
			7'd76: begin
				__main___storak76 <= convert_sync_array_muxed1;
			end
			7'd77: begin
				__main___storak77 <= convert_sync_array_muxed1;
			end
			7'd78: begin
				__main___storak78 <= convert_sync_array_muxed1;
			end
			7'd79: begin
				__main___storak79 <= convert_sync_array_muxed1;
			end
			7'd80: begin
				__main___storak80 <= convert_sync_array_muxed1;
			end
			7'd81: begin
				__main___storak81 <= convert_sync_array_muxed1;
			end
			7'd82: begin
				__main___storak82 <= convert_sync_array_muxed1;
			end
			7'd83: begin
				__main___storak83 <= convert_sync_array_muxed1;
			end
			7'd84: begin
				__main___storak84 <= convert_sync_array_muxed1;
			end
			7'd85: begin
				__main___storak85 <= convert_sync_array_muxed1;
			end
			7'd86: begin
				__main___storak86 <= convert_sync_array_muxed1;
			end
			7'd87: begin
				__main___storak87 <= convert_sync_array_muxed1;
			end
			7'd88: begin
				__main___storak88 <= convert_sync_array_muxed1;
			end
			7'd89: begin
				__main___storak89 <= convert_sync_array_muxed1;
			end
			7'd90: begin
				__main___storak90 <= convert_sync_array_muxed1;
			end
			7'd91: begin
				__main___storak91 <= convert_sync_array_muxed1;
			end
			7'd92: begin
				__main___storak92 <= convert_sync_array_muxed1;
			end
			7'd93: begin
				__main___storak93 <= convert_sync_array_muxed1;
			end
			7'd94: begin
				__main___storak94 <= convert_sync_array_muxed1;
			end
			7'd95: begin
				__main___storak95 <= convert_sync_array_muxed1;
			end
			7'd96: begin
				__main___storak96 <= convert_sync_array_muxed1;
			end
			7'd97: begin
				__main___storak97 <= convert_sync_array_muxed1;
			end
			7'd98: begin
				__main___storak98 <= convert_sync_array_muxed1;
			end
			7'd99: begin
				__main___storak99 <= convert_sync_array_muxed1;
			end
			7'd100: begin
				__main___storak100 <= convert_sync_array_muxed1;
			end
			7'd101: begin
				__main___storak101 <= convert_sync_array_muxed1;
			end
			7'd102: begin
				__main___storak102 <= convert_sync_array_muxed1;
			end
			7'd103: begin
				__main___storak103 <= convert_sync_array_muxed1;
			end
			7'd104: begin
				__main___storak104 <= convert_sync_array_muxed1;
			end
			7'd105: begin
				__main___storak105 <= convert_sync_array_muxed1;
			end
			7'd106: begin
				__main___storak106 <= convert_sync_array_muxed1;
			end
			7'd107: begin
				__main___storak107 <= convert_sync_array_muxed1;
			end
			7'd108: begin
				__main___storak108 <= convert_sync_array_muxed1;
			end
			7'd109: begin
				__main___storak109 <= convert_sync_array_muxed1;
			end
			7'd110: begin
				__main___storak110 <= convert_sync_array_muxed1;
			end
			7'd111: begin
				__main___storak111 <= convert_sync_array_muxed1;
			end
			7'd112: begin
				__main___storak112 <= convert_sync_array_muxed1;
			end
			7'd113: begin
				__main___storak113 <= convert_sync_array_muxed1;
			end
			7'd114: begin
				__main___storak114 <= convert_sync_array_muxed1;
			end
			7'd115: begin
				__main___storak115 <= convert_sync_array_muxed1;
			end
			7'd116: begin
				__main___storak116 <= convert_sync_array_muxed1;
			end
			7'd117: begin
				__main___storak117 <= convert_sync_array_muxed1;
			end
			7'd118: begin
				__main___storak118 <= convert_sync_array_muxed1;
			end
			7'd119: begin
				__main___storak119 <= convert_sync_array_muxed1;
			end
			7'd120: begin
				__main___storak120 <= convert_sync_array_muxed1;
			end
			7'd121: begin
				__main___storak121 <= convert_sync_array_muxed1;
			end
			7'd122: begin
				__main___storak122 <= convert_sync_array_muxed1;
			end
			7'd123: begin
				__main___storak123 <= convert_sync_array_muxed1;
			end
			7'd124: begin
				__main___storak124 <= convert_sync_array_muxed1;
			end
			7'd125: begin
				__main___storak125 <= convert_sync_array_muxed1;
			end
			7'd126: begin
				__main___storak126 <= convert_sync_array_muxed1;
			end
			default: begin
				__main___storak127 <= convert_sync_array_muxed1;
			end
		endcase
	end
	if (convert_t_next_value_ce) begin
		convert_sync_array_muxed2 = convert_t_next_value;
		case (ADR_i)
			1'd0: begin
				__main___storak0 <= convert_sync_array_muxed2;
			end
			1'd1: begin
				__main___storak1 <= convert_sync_array_muxed2;
			end
			2'd2: begin
				__main___storak2 <= convert_sync_array_muxed2;
			end
			2'd3: begin
				__main___storak3 <= convert_sync_array_muxed2;
			end
			3'd4: begin
				__main___storak4 <= convert_sync_array_muxed2;
			end
			3'd5: begin
				__main___storak5 <= convert_sync_array_muxed2;
			end
			3'd6: begin
				__main___storak6 <= convert_sync_array_muxed2;
			end
			3'd7: begin
				__main___storak7 <= convert_sync_array_muxed2;
			end
			4'd8: begin
				__main___storak8 <= convert_sync_array_muxed2;
			end
			4'd9: begin
				__main___storak9 <= convert_sync_array_muxed2;
			end
			4'd10: begin
				__main___storak10 <= convert_sync_array_muxed2;
			end
			4'd11: begin
				__main___storak11 <= convert_sync_array_muxed2;
			end
			4'd12: begin
				__main___storak12 <= convert_sync_array_muxed2;
			end
			4'd13: begin
				__main___storak13 <= convert_sync_array_muxed2;
			end
			4'd14: begin
				__main___storak14 <= convert_sync_array_muxed2;
			end
			4'd15: begin
				__main___storak15 <= convert_sync_array_muxed2;
			end
			5'd16: begin
				__main___storak16 <= convert_sync_array_muxed2;
			end
			5'd17: begin
				__main___storak17 <= convert_sync_array_muxed2;
			end
			5'd18: begin
				__main___storak18 <= convert_sync_array_muxed2;
			end
			5'd19: begin
				__main___storak19 <= convert_sync_array_muxed2;
			end
			5'd20: begin
				__main___storak20 <= convert_sync_array_muxed2;
			end
			5'd21: begin
				__main___storak21 <= convert_sync_array_muxed2;
			end
			5'd22: begin
				__main___storak22 <= convert_sync_array_muxed2;
			end
			5'd23: begin
				__main___storak23 <= convert_sync_array_muxed2;
			end
			5'd24: begin
				__main___storak24 <= convert_sync_array_muxed2;
			end
			5'd25: begin
				__main___storak25 <= convert_sync_array_muxed2;
			end
			5'd26: begin
				__main___storak26 <= convert_sync_array_muxed2;
			end
			5'd27: begin
				__main___storak27 <= convert_sync_array_muxed2;
			end
			5'd28: begin
				__main___storak28 <= convert_sync_array_muxed2;
			end
			5'd29: begin
				__main___storak29 <= convert_sync_array_muxed2;
			end
			5'd30: begin
				__main___storak30 <= convert_sync_array_muxed2;
			end
			5'd31: begin
				__main___storak31 <= convert_sync_array_muxed2;
			end
			6'd32: begin
				__main___storak32 <= convert_sync_array_muxed2;
			end
			6'd33: begin
				__main___storak33 <= convert_sync_array_muxed2;
			end
			6'd34: begin
				__main___storak34 <= convert_sync_array_muxed2;
			end
			6'd35: begin
				__main___storak35 <= convert_sync_array_muxed2;
			end
			6'd36: begin
				__main___storak36 <= convert_sync_array_muxed2;
			end
			6'd37: begin
				__main___storak37 <= convert_sync_array_muxed2;
			end
			6'd38: begin
				__main___storak38 <= convert_sync_array_muxed2;
			end
			6'd39: begin
				__main___storak39 <= convert_sync_array_muxed2;
			end
			6'd40: begin
				__main___storak40 <= convert_sync_array_muxed2;
			end
			6'd41: begin
				__main___storak41 <= convert_sync_array_muxed2;
			end
			6'd42: begin
				__main___storak42 <= convert_sync_array_muxed2;
			end
			6'd43: begin
				__main___storak43 <= convert_sync_array_muxed2;
			end
			6'd44: begin
				__main___storak44 <= convert_sync_array_muxed2;
			end
			6'd45: begin
				__main___storak45 <= convert_sync_array_muxed2;
			end
			6'd46: begin
				__main___storak46 <= convert_sync_array_muxed2;
			end
			6'd47: begin
				__main___storak47 <= convert_sync_array_muxed2;
			end
			6'd48: begin
				__main___storak48 <= convert_sync_array_muxed2;
			end
			6'd49: begin
				__main___storak49 <= convert_sync_array_muxed2;
			end
			6'd50: begin
				__main___storak50 <= convert_sync_array_muxed2;
			end
			6'd51: begin
				__main___storak51 <= convert_sync_array_muxed2;
			end
			6'd52: begin
				__main___storak52 <= convert_sync_array_muxed2;
			end
			6'd53: begin
				__main___storak53 <= convert_sync_array_muxed2;
			end
			6'd54: begin
				__main___storak54 <= convert_sync_array_muxed2;
			end
			6'd55: begin
				__main___storak55 <= convert_sync_array_muxed2;
			end
			6'd56: begin
				__main___storak56 <= convert_sync_array_muxed2;
			end
			6'd57: begin
				__main___storak57 <= convert_sync_array_muxed2;
			end
			6'd58: begin
				__main___storak58 <= convert_sync_array_muxed2;
			end
			6'd59: begin
				__main___storak59 <= convert_sync_array_muxed2;
			end
			6'd60: begin
				__main___storak60 <= convert_sync_array_muxed2;
			end
			6'd61: begin
				__main___storak61 <= convert_sync_array_muxed2;
			end
			6'd62: begin
				__main___storak62 <= convert_sync_array_muxed2;
			end
			6'd63: begin
				__main___storak63 <= convert_sync_array_muxed2;
			end
			7'd64: begin
				__main___storak64 <= convert_sync_array_muxed2;
			end
			7'd65: begin
				__main___storak65 <= convert_sync_array_muxed2;
			end
			7'd66: begin
				__main___storak66 <= convert_sync_array_muxed2;
			end
			7'd67: begin
				__main___storak67 <= convert_sync_array_muxed2;
			end
			7'd68: begin
				__main___storak68 <= convert_sync_array_muxed2;
			end
			7'd69: begin
				__main___storak69 <= convert_sync_array_muxed2;
			end
			7'd70: begin
				__main___storak70 <= convert_sync_array_muxed2;
			end
			7'd71: begin
				__main___storak71 <= convert_sync_array_muxed2;
			end
			7'd72: begin
				__main___storak72 <= convert_sync_array_muxed2;
			end
			7'd73: begin
				__main___storak73 <= convert_sync_array_muxed2;
			end
			7'd74: begin
				__main___storak74 <= convert_sync_array_muxed2;
			end
			7'd75: begin
				__main___storak75 <= convert_sync_array_muxed2;
			end
			7'd76: begin
				__main___storak76 <= convert_sync_array_muxed2;
			end
			7'd77: begin
				__main___storak77 <= convert_sync_array_muxed2;
			end
			7'd78: begin
				__main___storak78 <= convert_sync_array_muxed2;
			end
			7'd79: begin
				__main___storak79 <= convert_sync_array_muxed2;
			end
			7'd80: begin
				__main___storak80 <= convert_sync_array_muxed2;
			end
			7'd81: begin
				__main___storak81 <= convert_sync_array_muxed2;
			end
			7'd82: begin
				__main___storak82 <= convert_sync_array_muxed2;
			end
			7'd83: begin
				__main___storak83 <= convert_sync_array_muxed2;
			end
			7'd84: begin
				__main___storak84 <= convert_sync_array_muxed2;
			end
			7'd85: begin
				__main___storak85 <= convert_sync_array_muxed2;
			end
			7'd86: begin
				__main___storak86 <= convert_sync_array_muxed2;
			end
			7'd87: begin
				__main___storak87 <= convert_sync_array_muxed2;
			end
			7'd88: begin
				__main___storak88 <= convert_sync_array_muxed2;
			end
			7'd89: begin
				__main___storak89 <= convert_sync_array_muxed2;
			end
			7'd90: begin
				__main___storak90 <= convert_sync_array_muxed2;
			end
			7'd91: begin
				__main___storak91 <= convert_sync_array_muxed2;
			end
			7'd92: begin
				__main___storak92 <= convert_sync_array_muxed2;
			end
			7'd93: begin
				__main___storak93 <= convert_sync_array_muxed2;
			end
			7'd94: begin
				__main___storak94 <= convert_sync_array_muxed2;
			end
			7'd95: begin
				__main___storak95 <= convert_sync_array_muxed2;
			end
			7'd96: begin
				__main___storak96 <= convert_sync_array_muxed2;
			end
			7'd97: begin
				__main___storak97 <= convert_sync_array_muxed2;
			end
			7'd98: begin
				__main___storak98 <= convert_sync_array_muxed2;
			end
			7'd99: begin
				__main___storak99 <= convert_sync_array_muxed2;
			end
			7'd100: begin
				__main___storak100 <= convert_sync_array_muxed2;
			end
			7'd101: begin
				__main___storak101 <= convert_sync_array_muxed2;
			end
			7'd102: begin
				__main___storak102 <= convert_sync_array_muxed2;
			end
			7'd103: begin
				__main___storak103 <= convert_sync_array_muxed2;
			end
			7'd104: begin
				__main___storak104 <= convert_sync_array_muxed2;
			end
			7'd105: begin
				__main___storak105 <= convert_sync_array_muxed2;
			end
			7'd106: begin
				__main___storak106 <= convert_sync_array_muxed2;
			end
			7'd107: begin
				__main___storak107 <= convert_sync_array_muxed2;
			end
			7'd108: begin
				__main___storak108 <= convert_sync_array_muxed2;
			end
			7'd109: begin
				__main___storak109 <= convert_sync_array_muxed2;
			end
			7'd110: begin
				__main___storak110 <= convert_sync_array_muxed2;
			end
			7'd111: begin
				__main___storak111 <= convert_sync_array_muxed2;
			end
			7'd112: begin
				__main___storak112 <= convert_sync_array_muxed2;
			end
			7'd113: begin
				__main___storak113 <= convert_sync_array_muxed2;
			end
			7'd114: begin
				__main___storak114 <= convert_sync_array_muxed2;
			end
			7'd115: begin
				__main___storak115 <= convert_sync_array_muxed2;
			end
			7'd116: begin
				__main___storak116 <= convert_sync_array_muxed2;
			end
			7'd117: begin
				__main___storak117 <= convert_sync_array_muxed2;
			end
			7'd118: begin
				__main___storak118 <= convert_sync_array_muxed2;
			end
			7'd119: begin
				__main___storak119 <= convert_sync_array_muxed2;
			end
			7'd120: begin
				__main___storak120 <= convert_sync_array_muxed2;
			end
			7'd121: begin
				__main___storak121 <= convert_sync_array_muxed2;
			end
			7'd122: begin
				__main___storak122 <= convert_sync_array_muxed2;
			end
			7'd123: begin
				__main___storak123 <= convert_sync_array_muxed2;
			end
			7'd124: begin
				__main___storak124 <= convert_sync_array_muxed2;
			end
			7'd125: begin
				__main___storak125 <= convert_sync_array_muxed2;
			end
			7'd126: begin
				__main___storak126 <= convert_sync_array_muxed2;
			end
			default: begin
				__main___storak127 <= convert_sync_array_muxed2;
			end
		endcase
	end
	if (convert_f_next_value_ce) begin
		convert_sync_array_muxed3 = convert_f_next_value;
		case (ADR_i)
			1'd0: begin
				__main___storav0 <= convert_sync_array_muxed3;
			end
			1'd1: begin
				__main___storav1 <= convert_sync_array_muxed3;
			end
			2'd2: begin
				__main___storav2 <= convert_sync_array_muxed3;
			end
			2'd3: begin
				__main___storav3 <= convert_sync_array_muxed3;
			end
			3'd4: begin
				__main___storav4 <= convert_sync_array_muxed3;
			end
			3'd5: begin
				__main___storav5 <= convert_sync_array_muxed3;
			end
			3'd6: begin
				__main___storav6 <= convert_sync_array_muxed3;
			end
			3'd7: begin
				__main___storav7 <= convert_sync_array_muxed3;
			end
			4'd8: begin
				__main___storav8 <= convert_sync_array_muxed3;
			end
			4'd9: begin
				__main___storav9 <= convert_sync_array_muxed3;
			end
			4'd10: begin
				__main___storav10 <= convert_sync_array_muxed3;
			end
			4'd11: begin
				__main___storav11 <= convert_sync_array_muxed3;
			end
			4'd12: begin
				__main___storav12 <= convert_sync_array_muxed3;
			end
			4'd13: begin
				__main___storav13 <= convert_sync_array_muxed3;
			end
			4'd14: begin
				__main___storav14 <= convert_sync_array_muxed3;
			end
			4'd15: begin
				__main___storav15 <= convert_sync_array_muxed3;
			end
			5'd16: begin
				__main___storav16 <= convert_sync_array_muxed3;
			end
			5'd17: begin
				__main___storav17 <= convert_sync_array_muxed3;
			end
			5'd18: begin
				__main___storav18 <= convert_sync_array_muxed3;
			end
			5'd19: begin
				__main___storav19 <= convert_sync_array_muxed3;
			end
			5'd20: begin
				__main___storav20 <= convert_sync_array_muxed3;
			end
			5'd21: begin
				__main___storav21 <= convert_sync_array_muxed3;
			end
			5'd22: begin
				__main___storav22 <= convert_sync_array_muxed3;
			end
			5'd23: begin
				__main___storav23 <= convert_sync_array_muxed3;
			end
			5'd24: begin
				__main___storav24 <= convert_sync_array_muxed3;
			end
			5'd25: begin
				__main___storav25 <= convert_sync_array_muxed3;
			end
			5'd26: begin
				__main___storav26 <= convert_sync_array_muxed3;
			end
			5'd27: begin
				__main___storav27 <= convert_sync_array_muxed3;
			end
			5'd28: begin
				__main___storav28 <= convert_sync_array_muxed3;
			end
			5'd29: begin
				__main___storav29 <= convert_sync_array_muxed3;
			end
			5'd30: begin
				__main___storav30 <= convert_sync_array_muxed3;
			end
			5'd31: begin
				__main___storav31 <= convert_sync_array_muxed3;
			end
			6'd32: begin
				__main___storav32 <= convert_sync_array_muxed3;
			end
			6'd33: begin
				__main___storav33 <= convert_sync_array_muxed3;
			end
			6'd34: begin
				__main___storav34 <= convert_sync_array_muxed3;
			end
			6'd35: begin
				__main___storav35 <= convert_sync_array_muxed3;
			end
			6'd36: begin
				__main___storav36 <= convert_sync_array_muxed3;
			end
			6'd37: begin
				__main___storav37 <= convert_sync_array_muxed3;
			end
			6'd38: begin
				__main___storav38 <= convert_sync_array_muxed3;
			end
			6'd39: begin
				__main___storav39 <= convert_sync_array_muxed3;
			end
			6'd40: begin
				__main___storav40 <= convert_sync_array_muxed3;
			end
			6'd41: begin
				__main___storav41 <= convert_sync_array_muxed3;
			end
			6'd42: begin
				__main___storav42 <= convert_sync_array_muxed3;
			end
			6'd43: begin
				__main___storav43 <= convert_sync_array_muxed3;
			end
			6'd44: begin
				__main___storav44 <= convert_sync_array_muxed3;
			end
			6'd45: begin
				__main___storav45 <= convert_sync_array_muxed3;
			end
			6'd46: begin
				__main___storav46 <= convert_sync_array_muxed3;
			end
			6'd47: begin
				__main___storav47 <= convert_sync_array_muxed3;
			end
			6'd48: begin
				__main___storav48 <= convert_sync_array_muxed3;
			end
			6'd49: begin
				__main___storav49 <= convert_sync_array_muxed3;
			end
			6'd50: begin
				__main___storav50 <= convert_sync_array_muxed3;
			end
			6'd51: begin
				__main___storav51 <= convert_sync_array_muxed3;
			end
			6'd52: begin
				__main___storav52 <= convert_sync_array_muxed3;
			end
			6'd53: begin
				__main___storav53 <= convert_sync_array_muxed3;
			end
			6'd54: begin
				__main___storav54 <= convert_sync_array_muxed3;
			end
			6'd55: begin
				__main___storav55 <= convert_sync_array_muxed3;
			end
			6'd56: begin
				__main___storav56 <= convert_sync_array_muxed3;
			end
			6'd57: begin
				__main___storav57 <= convert_sync_array_muxed3;
			end
			6'd58: begin
				__main___storav58 <= convert_sync_array_muxed3;
			end
			6'd59: begin
				__main___storav59 <= convert_sync_array_muxed3;
			end
			6'd60: begin
				__main___storav60 <= convert_sync_array_muxed3;
			end
			6'd61: begin
				__main___storav61 <= convert_sync_array_muxed3;
			end
			6'd62: begin
				__main___storav62 <= convert_sync_array_muxed3;
			end
			6'd63: begin
				__main___storav63 <= convert_sync_array_muxed3;
			end
			7'd64: begin
				__main___storav64 <= convert_sync_array_muxed3;
			end
			7'd65: begin
				__main___storav65 <= convert_sync_array_muxed3;
			end
			7'd66: begin
				__main___storav66 <= convert_sync_array_muxed3;
			end
			7'd67: begin
				__main___storav67 <= convert_sync_array_muxed3;
			end
			7'd68: begin
				__main___storav68 <= convert_sync_array_muxed3;
			end
			7'd69: begin
				__main___storav69 <= convert_sync_array_muxed3;
			end
			7'd70: begin
				__main___storav70 <= convert_sync_array_muxed3;
			end
			7'd71: begin
				__main___storav71 <= convert_sync_array_muxed3;
			end
			7'd72: begin
				__main___storav72 <= convert_sync_array_muxed3;
			end
			7'd73: begin
				__main___storav73 <= convert_sync_array_muxed3;
			end
			7'd74: begin
				__main___storav74 <= convert_sync_array_muxed3;
			end
			7'd75: begin
				__main___storav75 <= convert_sync_array_muxed3;
			end
			7'd76: begin
				__main___storav76 <= convert_sync_array_muxed3;
			end
			7'd77: begin
				__main___storav77 <= convert_sync_array_muxed3;
			end
			7'd78: begin
				__main___storav78 <= convert_sync_array_muxed3;
			end
			7'd79: begin
				__main___storav79 <= convert_sync_array_muxed3;
			end
			7'd80: begin
				__main___storav80 <= convert_sync_array_muxed3;
			end
			7'd81: begin
				__main___storav81 <= convert_sync_array_muxed3;
			end
			7'd82: begin
				__main___storav82 <= convert_sync_array_muxed3;
			end
			7'd83: begin
				__main___storav83 <= convert_sync_array_muxed3;
			end
			7'd84: begin
				__main___storav84 <= convert_sync_array_muxed3;
			end
			7'd85: begin
				__main___storav85 <= convert_sync_array_muxed3;
			end
			7'd86: begin
				__main___storav86 <= convert_sync_array_muxed3;
			end
			7'd87: begin
				__main___storav87 <= convert_sync_array_muxed3;
			end
			7'd88: begin
				__main___storav88 <= convert_sync_array_muxed3;
			end
			7'd89: begin
				__main___storav89 <= convert_sync_array_muxed3;
			end
			7'd90: begin
				__main___storav90 <= convert_sync_array_muxed3;
			end
			7'd91: begin
				__main___storav91 <= convert_sync_array_muxed3;
			end
			7'd92: begin
				__main___storav92 <= convert_sync_array_muxed3;
			end
			7'd93: begin
				__main___storav93 <= convert_sync_array_muxed3;
			end
			7'd94: begin
				__main___storav94 <= convert_sync_array_muxed3;
			end
			7'd95: begin
				__main___storav95 <= convert_sync_array_muxed3;
			end
			7'd96: begin
				__main___storav96 <= convert_sync_array_muxed3;
			end
			7'd97: begin
				__main___storav97 <= convert_sync_array_muxed3;
			end
			7'd98: begin
				__main___storav98 <= convert_sync_array_muxed3;
			end
			7'd99: begin
				__main___storav99 <= convert_sync_array_muxed3;
			end
			7'd100: begin
				__main___storav100 <= convert_sync_array_muxed3;
			end
			7'd101: begin
				__main___storav101 <= convert_sync_array_muxed3;
			end
			7'd102: begin
				__main___storav102 <= convert_sync_array_muxed3;
			end
			7'd103: begin
				__main___storav103 <= convert_sync_array_muxed3;
			end
			7'd104: begin
				__main___storav104 <= convert_sync_array_muxed3;
			end
			7'd105: begin
				__main___storav105 <= convert_sync_array_muxed3;
			end
			7'd106: begin
				__main___storav106 <= convert_sync_array_muxed3;
			end
			7'd107: begin
				__main___storav107 <= convert_sync_array_muxed3;
			end
			7'd108: begin
				__main___storav108 <= convert_sync_array_muxed3;
			end
			7'd109: begin
				__main___storav109 <= convert_sync_array_muxed3;
			end
			7'd110: begin
				__main___storav110 <= convert_sync_array_muxed3;
			end
			7'd111: begin
				__main___storav111 <= convert_sync_array_muxed3;
			end
			7'd112: begin
				__main___storav112 <= convert_sync_array_muxed3;
			end
			7'd113: begin
				__main___storav113 <= convert_sync_array_muxed3;
			end
			7'd114: begin
				__main___storav114 <= convert_sync_array_muxed3;
			end
			7'd115: begin
				__main___storav115 <= convert_sync_array_muxed3;
			end
			7'd116: begin
				__main___storav116 <= convert_sync_array_muxed3;
			end
			7'd117: begin
				__main___storav117 <= convert_sync_array_muxed3;
			end
			7'd118: begin
				__main___storav118 <= convert_sync_array_muxed3;
			end
			7'd119: begin
				__main___storav119 <= convert_sync_array_muxed3;
			end
			7'd120: begin
				__main___storav120 <= convert_sync_array_muxed3;
			end
			7'd121: begin
				__main___storav121 <= convert_sync_array_muxed3;
			end
			7'd122: begin
				__main___storav122 <= convert_sync_array_muxed3;
			end
			7'd123: begin
				__main___storav123 <= convert_sync_array_muxed3;
			end
			7'd124: begin
				__main___storav124 <= convert_sync_array_muxed3;
			end
			7'd125: begin
				__main___storav125 <= convert_sync_array_muxed3;
			end
			7'd126: begin
				__main___storav126 <= convert_sync_array_muxed3;
			end
			default: begin
				__main___storav127 <= convert_sync_array_muxed3;
			end
		endcase
	end
	if (sys_rst_1) begin
		STALL_o <= 1'd0;
		ACK_o <= 1'd0;
		DAT_o <= 64'd0;
		__main___storak0 <= 64'd0;
		__main___storak1 <= 64'd0;
		__main___storak2 <= 64'd0;
		__main___storak3 <= 64'd0;
		__main___storak4 <= 64'd0;
		__main___storak5 <= 64'd0;
		__main___storak6 <= 64'd0;
		__main___storak7 <= 64'd0;
		__main___storak8 <= 64'd0;
		__main___storak9 <= 64'd0;
		__main___storak10 <= 64'd0;
		__main___storak11 <= 64'd0;
		__main___storak12 <= 64'd0;
		__main___storak13 <= 64'd0;
		__main___storak14 <= 64'd0;
		__main___storak15 <= 64'd0;
		__main___storak16 <= 64'd0;
		__main___storak17 <= 64'd0;
		__main___storak18 <= 64'd0;
		__main___storak19 <= 64'd0;
		__main___storak20 <= 64'd0;
		__main___storak21 <= 64'd0;
		__main___storak22 <= 64'd0;
		__main___storak23 <= 64'd0;
		__main___storak24 <= 64'd0;
		__main___storak25 <= 64'd0;
		__main___storak26 <= 64'd0;
		__main___storak27 <= 64'd0;
		__main___storak28 <= 64'd0;
		__main___storak29 <= 64'd0;
		__main___storak30 <= 64'd0;
		__main___storak31 <= 64'd0;
		__main___storak32 <= 64'd0;
		__main___storak33 <= 64'd0;
		__main___storak34 <= 64'd0;
		__main___storak35 <= 64'd0;
		__main___storak36 <= 64'd0;
		__main___storak37 <= 64'd0;
		__main___storak38 <= 64'd0;
		__main___storak39 <= 64'd0;
		__main___storak40 <= 64'd0;
		__main___storak41 <= 64'd0;
		__main___storak42 <= 64'd0;
		__main___storak43 <= 64'd0;
		__main___storak44 <= 64'd0;
		__main___storak45 <= 64'd0;
		__main___storak46 <= 64'd0;
		__main___storak47 <= 64'd0;
		__main___storak48 <= 64'd0;
		__main___storak49 <= 64'd0;
		__main___storak50 <= 64'd0;
		__main___storak51 <= 64'd0;
		__main___storak52 <= 64'd0;
		__main___storak53 <= 64'd0;
		__main___storak54 <= 64'd0;
		__main___storak55 <= 64'd0;
		__main___storak56 <= 64'd0;
		__main___storak57 <= 64'd0;
		__main___storak58 <= 64'd0;
		__main___storak59 <= 64'd0;
		__main___storak60 <= 64'd0;
		__main___storak61 <= 64'd0;
		__main___storak62 <= 64'd0;
		__main___storak63 <= 64'd0;
		__main___storak64 <= 64'd0;
		__main___storak65 <= 64'd0;
		__main___storak66 <= 64'd0;
		__main___storak67 <= 64'd0;
		__main___storak68 <= 64'd0;
		__main___storak69 <= 64'd0;
		__main___storak70 <= 64'd0;
		__main___storak71 <= 64'd0;
		__main___storak72 <= 64'd0;
		__main___storak73 <= 64'd0;
		__main___storak74 <= 64'd0;
		__main___storak75 <= 64'd0;
		__main___storak76 <= 64'd0;
		__main___storak77 <= 64'd0;
		__main___storak78 <= 64'd0;
		__main___storak79 <= 64'd0;
		__main___storak80 <= 64'd0;
		__main___storak81 <= 64'd0;
		__main___storak82 <= 64'd0;
		__main___storak83 <= 64'd0;
		__main___storak84 <= 64'd0;
		__main___storak85 <= 64'd0;
		__main___storak86 <= 64'd0;
		__main___storak87 <= 64'd0;
		__main___storak88 <= 64'd0;
		__main___storak89 <= 64'd0;
		__main___storak90 <= 64'd0;
		__main___storak91 <= 64'd0;
		__main___storak92 <= 64'd0;
		__main___storak93 <= 64'd0;
		__main___storak94 <= 64'd0;
		__main___storak95 <= 64'd0;
		__main___storak96 <= 64'd0;
		__main___storak97 <= 64'd0;
		__main___storak98 <= 64'd0;
		__main___storak99 <= 64'd0;
		__main___storak100 <= 64'd0;
		__main___storak101 <= 64'd0;
		__main___storak102 <= 64'd0;
		__main___storak103 <= 64'd0;
		__main___storak104 <= 64'd0;
		__main___storak105 <= 64'd0;
		__main___storak106 <= 64'd0;
		__main___storak107 <= 64'd0;
		__main___storak108 <= 64'd0;
		__main___storak109 <= 64'd0;
		__main___storak110 <= 64'd0;
		__main___storak111 <= 64'd0;
		__main___storak112 <= 64'd0;
		__main___storak113 <= 64'd0;
		__main___storak114 <= 64'd0;
		__main___storak115 <= 64'd0;
		__main___storak116 <= 64'd0;
		__main___storak117 <= 64'd0;
		__main___storak118 <= 64'd0;
		__main___storak119 <= 64'd0;
		__main___storak120 <= 64'd0;
		__main___storak121 <= 64'd0;
		__main___storak122 <= 64'd0;
		__main___storak123 <= 64'd0;
		__main___storak124 <= 64'd0;
		__main___storak125 <= 64'd0;
		__main___storak126 <= 64'd0;
		__main___storak127 <= 64'd0;
		__main___storav0 <= 64'd0;
		__main___storav1 <= 64'd0;
		__main___storav2 <= 64'd0;
		__main___storav3 <= 64'd0;
		__main___storav4 <= 64'd0;
		__main___storav5 <= 64'd0;
		__main___storav6 <= 64'd0;
		__main___storav7 <= 64'd0;
		__main___storav8 <= 64'd0;
		__main___storav9 <= 64'd0;
		__main___storav10 <= 64'd0;
		__main___storav11 <= 64'd0;
		__main___storav12 <= 64'd0;
		__main___storav13 <= 64'd0;
		__main___storav14 <= 64'd0;
		__main___storav15 <= 64'd0;
		__main___storav16 <= 64'd0;
		__main___storav17 <= 64'd0;
		__main___storav18 <= 64'd0;
		__main___storav19 <= 64'd0;
		__main___storav20 <= 64'd0;
		__main___storav21 <= 64'd0;
		__main___storav22 <= 64'd0;
		__main___storav23 <= 64'd0;
		__main___storav24 <= 64'd0;
		__main___storav25 <= 64'd0;
		__main___storav26 <= 64'd0;
		__main___storav27 <= 64'd0;
		__main___storav28 <= 64'd0;
		__main___storav29 <= 64'd0;
		__main___storav30 <= 64'd0;
		__main___storav31 <= 64'd0;
		__main___storav32 <= 64'd0;
		__main___storav33 <= 64'd0;
		__main___storav34 <= 64'd0;
		__main___storav35 <= 64'd0;
		__main___storav36 <= 64'd0;
		__main___storav37 <= 64'd0;
		__main___storav38 <= 64'd0;
		__main___storav39 <= 64'd0;
		__main___storav40 <= 64'd0;
		__main___storav41 <= 64'd0;
		__main___storav42 <= 64'd0;
		__main___storav43 <= 64'd0;
		__main___storav44 <= 64'd0;
		__main___storav45 <= 64'd0;
		__main___storav46 <= 64'd0;
		__main___storav47 <= 64'd0;
		__main___storav48 <= 64'd0;
		__main___storav49 <= 64'd0;
		__main___storav50 <= 64'd0;
		__main___storav51 <= 64'd0;
		__main___storav52 <= 64'd0;
		__main___storav53 <= 64'd0;
		__main___storav54 <= 64'd0;
		__main___storav55 <= 64'd0;
		__main___storav56 <= 64'd0;
		__main___storav57 <= 64'd0;
		__main___storav58 <= 64'd0;
		__main___storav59 <= 64'd0;
		__main___storav60 <= 64'd0;
		__main___storav61 <= 64'd0;
		__main___storav62 <= 64'd0;
		__main___storav63 <= 64'd0;
		__main___storav64 <= 64'd0;
		__main___storav65 <= 64'd0;
		__main___storav66 <= 64'd0;
		__main___storav67 <= 64'd0;
		__main___storav68 <= 64'd0;
		__main___storav69 <= 64'd0;
		__main___storav70 <= 64'd0;
		__main___storav71 <= 64'd0;
		__main___storav72 <= 64'd0;
		__main___storav73 <= 64'd0;
		__main___storav74 <= 64'd0;
		__main___storav75 <= 64'd0;
		__main___storav76 <= 64'd0;
		__main___storav77 <= 64'd0;
		__main___storav78 <= 64'd0;
		__main___storav79 <= 64'd0;
		__main___storav80 <= 64'd0;
		__main___storav81 <= 64'd0;
		__main___storav82 <= 64'd0;
		__main___storav83 <= 64'd0;
		__main___storav84 <= 64'd0;
		__main___storav85 <= 64'd0;
		__main___storav86 <= 64'd0;
		__main___storav87 <= 64'd0;
		__main___storav88 <= 64'd0;
		__main___storav89 <= 64'd0;
		__main___storav90 <= 64'd0;
		__main___storav91 <= 64'd0;
		__main___storav92 <= 64'd0;
		__main___storav93 <= 64'd0;
		__main___storav94 <= 64'd0;
		__main___storav95 <= 64'd0;
		__main___storav96 <= 64'd0;
		__main___storav97 <= 64'd0;
		__main___storav98 <= 64'd0;
		__main___storav99 <= 64'd0;
		__main___storav100 <= 64'd0;
		__main___storav101 <= 64'd0;
		__main___storav102 <= 64'd0;
		__main___storav103 <= 64'd0;
		__main___storav104 <= 64'd0;
		__main___storav105 <= 64'd0;
		__main___storav106 <= 64'd0;
		__main___storav107 <= 64'd0;
		__main___storav108 <= 64'd0;
		__main___storav109 <= 64'd0;
		__main___storav110 <= 64'd0;
		__main___storav111 <= 64'd0;
		__main___storav112 <= 64'd0;
		__main___storav113 <= 64'd0;
		__main___storav114 <= 64'd0;
		__main___storav115 <= 64'd0;
		__main___storav116 <= 64'd0;
		__main___storav117 <= 64'd0;
		__main___storav118 <= 64'd0;
		__main___storav119 <= 64'd0;
		__main___storav120 <= 64'd0;
		__main___storav121 <= 64'd0;
		__main___storav122 <= 64'd0;
		__main___storav123 <= 64'd0;
		__main___storav124 <= 64'd0;
		__main___storav125 <= 64'd0;
		__main___storav126 <= 64'd0;
		__main___storav127 <= 64'd0;
		__main___empty_location <= 64'd0;
		convert_state <= 2'd3;
	end
end

endmodule


